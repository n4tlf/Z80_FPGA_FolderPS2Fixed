// Copyright (C) 2021  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 21.1.0 Build 842 10/21/2021 SJ Lite Edition"
// CREATED		"Wed Mar 30 13:44:51 2022"

module Z80_FPGA(
	CLK_50,
	FPGA_IN_XRDY,
	FPGA_IN_RDY,
	FPGA_IN_SDSB-,
	FPGA_IN_CDSB-,
	FPGA_IN_pHOLD-,
	FPGA_IN_DI0,
	FPGA_IN_DI1,
	FPGA_IN_DI2,
	FPGA_IN_DI4,
	FPGA_IN_DI5,
	FPGA_IN_DI6,
	FPGA_IN_DI7,
	FPGA_IN_DI3,
	FPGA_IN_PS2_CLK,
	FPGA_IN_PS2_DATA,
	FPGA_IN_PRN_ACK,
	FPGA_IN_PRN_BUSY,
	RTC_SPI_SO,
	DIP7,
	DIP6,
	DIP5,
	DIP4,
	DIP3,
	DIP2,
	DIP1,
	DIP0,
	FPGA_IN_INT_B-,
	FPGA_IN_INT_C-,
	FPGA_IN_INT_D-,
	FPGA_IN_INT_A-,
	USB_RX,
	FPGA_IN_INT-,
	RTC_INT,
	FPGA_IN_ENABLE_INTA,
	FPGA_IN_BOARD_RESET-,
	SD_DO,
	FPGA_OUT_A1,
	FPGA_OUT_A2,
	FPGA_OUT_A3,
	FPGA_OUT_A4,
	FPGA_OUT_A5,
	FPGA_OUT_A6,
	FPGA_OUT_A7,
	FPGA_OUT_A16,
	FPGA_OUT_A17,
	FPGA_OUT_A18,
	FPGA_OUT_A19,
	FPGA_OUT_CPU_CLK,
	FPGA_OUT_sINTA,
	FPGA_OUT_sM1,
	FPGA_OUT_sWO-,
	FPGA_OUT_sMEMR,
	FPGA_OUT_sINP,
	FPGA_OUT_sOUT,
	FPGA_OUT_sHLTA,
	FPGA_OUT_pDBIN,
	FPGA_OUT_pWR-,
	FPGA_OUT_MWRT,
	FPGA_OUT_2mHz_CLOCK,
	FPGA_OUT_PHI,
	FPGA_OUT_pSYNC,
	FPGA_OUT_pSTVAL-,
	FPGA_OUT_RAM_WR-,
	FPGA_OUT_RAM_OE-,
	FPGA_OUT_DO0,
	FPGA_OUT_DO1,
	FPGA_OUT_DO2,
	FPGA_OUT_DO3,
	FPGA_OUT_DO4,
	FPGA_OUT_DO5,
	FPGA_OUT_DO6,
	FPGA_OUT_DO7,
	FPGA_OUT_A0,
	FPGA_OUT_A8,
	FPGA_OUT_A9,
	FPGA_OUT_A11,
	FPGA_OUT_A10,
	FPGA_OUT_A12,
	FPGA_OUT_A13,
	FPGA_OUT_A14,
	FPGA_OUT_A15,
	FPGA_OUT_STATUS_DISABLE,
	FPGA_OUT_pHLDA,
	FPGA_OUT_CTL_DISABLE,
	FPGA_OUT_CTL_OE-,
	FPGA_OUT_STATUS_OE-,
	FPGA_ADD_OE-,
	FPGA_OUT_DO_OE-,
	FPGA_OUT_DI_OE-,
	FPGA_OUT_RAM_CS-,
	FPGA_OUT_RAM_A17,
	FPGA_OUT_RAM_A18,
	FPGA_OUT_RAM_A16,
	USB_TX,
	F_BAR0,
	F_BAR1,
	F_BAR2,
	F_BAR3,
	F_BAR4,
	F_BAR5,
	F_BAR6,
	F_BAR7,
	USB_TX_BUSY_LED,
	USB_RX_BUSY_LED,
	5V_OUT_IDE_PORTS_RD-,
	5V_OUT_IDE_PORTS_WR-,
	VGA_R,
	VGA_G,
	VGA_B,
	HSync,
	VSync,
	BUZZER,
	F_BOARD_ACTIVE-,
	FPGA_OUT_PRN_0,
	FPGA_OUT_PRN_1,
	FPGA_OUT_PRN_2,
	FPGA_OUT_PRN_3,
	FPGA_OUT_PRN_4,
	FPGA_OUT_PRN_5,
	FPGA_OUT_PRN_6,
	FPGA_OUT_PRN_7,
	FPGA_OUT_PRN_STROBE,
	PRN_ACK_LED,
	FPGA_OUT_PHANTOM,
	S100_PHANTOM_LED,
	RTC_CS,
	RTC_SPI_SI,
	RTC_SPI_CLK,
	SD_CMD,
	SD_CLK,
	LED_4,
	P1,
	LED_1,
	DIAG_LED,
	SD_CS_B-,
	FPGA_OUT_SPARE1,
	SD_CS_A-,
	FPGA_OUT_IDE_RD-,
	FPGA_OUT_IDE_WR-,
	FPGA_OUT_8255_SEL-,
	FPGA_OUT_HIGH_ROM_LED-,
	FPGA_OUT_LOW_ROM_LED-,
	FPGA_OUT_HIGH_RAM_LED-,
	LED_2,
	LED_3,
	FPGA_BI_D0,
	FPGA_BI_D1,
	FPGA_BI_D2,
	FPGA_BI_D3,
	FPGA_BI_D4,
	FPGA_BI_D5,
	FPGA_BI_D6,
	FPGA_BI_D7
);


input wire	CLK_50;
input wire	FPGA_IN_XRDY;
input wire	FPGA_IN_RDY;
input wire	FPGA_IN_SDSB-;
input wire	FPGA_IN_CDSB-;
input wire	FPGA_IN_pHOLD-;
input wire	FPGA_IN_DI0;
input wire	FPGA_IN_DI1;
input wire	FPGA_IN_DI2;
input wire	FPGA_IN_DI4;
input wire	FPGA_IN_DI5;
input wire	FPGA_IN_DI6;
input wire	FPGA_IN_DI7;
input wire	FPGA_IN_DI3;
input wire	FPGA_IN_PS2_CLK;
input wire	FPGA_IN_PS2_DATA;
input wire	FPGA_IN_PRN_ACK;
input wire	FPGA_IN_PRN_BUSY;
input wire	RTC_SPI_SO;
input wire	DIP7;
input wire	DIP6;
input wire	DIP5;
input wire	DIP4;
input wire	DIP3;
input wire	DIP2;
input wire	DIP1;
input wire	DIP0;
input wire	FPGA_IN_INT_B-;
input wire	FPGA_IN_INT_C-;
input wire	FPGA_IN_INT_D-;
input wire	FPGA_IN_INT_A-;
input wire	USB_RX;
input wire	FPGA_IN_INT-;
input wire	RTC_INT;
input wire	FPGA_IN_ENABLE_INTA;
input wire	FPGA_IN_BOARD_RESET-;
input wire	SD_DO;
output wire	FPGA_OUT_A1;
output wire	FPGA_OUT_A2;
output wire	FPGA_OUT_A3;
output wire	FPGA_OUT_A4;
output wire	FPGA_OUT_A5;
output wire	FPGA_OUT_A6;
output wire	FPGA_OUT_A7;
output wire	FPGA_OUT_A16;
output wire	FPGA_OUT_A17;
output wire	FPGA_OUT_A18;
output wire	FPGA_OUT_A19;
output wire	FPGA_OUT_CPU_CLK;
output wire	FPGA_OUT_sINTA;
output wire	FPGA_OUT_sM1;
output wire	FPGA_OUT_sWO-;
output wire	FPGA_OUT_sMEMR;
output wire	FPGA_OUT_sINP;
output wire	FPGA_OUT_sOUT;
output wire	FPGA_OUT_sHLTA;
output wire	FPGA_OUT_pDBIN;
output wire	FPGA_OUT_pWR-;
output wire	FPGA_OUT_MWRT;
output wire	FPGA_OUT_2mHz_CLOCK;
output wire	FPGA_OUT_PHI;
output wire	FPGA_OUT_pSYNC;
output wire	FPGA_OUT_pSTVAL-;
output wire	FPGA_OUT_RAM_WR-;
output wire	FPGA_OUT_RAM_OE-;
output wire	FPGA_OUT_DO0;
output wire	FPGA_OUT_DO1;
output wire	FPGA_OUT_DO2;
output wire	FPGA_OUT_DO3;
output wire	FPGA_OUT_DO4;
output wire	FPGA_OUT_DO5;
output wire	FPGA_OUT_DO6;
output wire	FPGA_OUT_DO7;
output wire	FPGA_OUT_A0;
output wire	FPGA_OUT_A8;
output wire	FPGA_OUT_A9;
output wire	FPGA_OUT_A11;
output wire	FPGA_OUT_A10;
output wire	FPGA_OUT_A12;
output wire	FPGA_OUT_A13;
output wire	FPGA_OUT_A14;
output wire	FPGA_OUT_A15;
output wire	FPGA_OUT_STATUS_DISABLE;
output wire	FPGA_OUT_pHLDA;
output wire	FPGA_OUT_CTL_DISABLE;
output wire	FPGA_OUT_CTL_OE-;
output wire	FPGA_OUT_STATUS_OE-;
output wire	FPGA_ADD_OE-;
output wire	FPGA_OUT_DO_OE-;
output wire	FPGA_OUT_DI_OE-;
output wire	FPGA_OUT_RAM_CS-;
output wire	FPGA_OUT_RAM_A17;
output wire	FPGA_OUT_RAM_A18;
output wire	FPGA_OUT_RAM_A16;
output wire	USB_TX;
output wire	F_BAR0;
output wire	F_BAR1;
output wire	F_BAR2;
output wire	F_BAR3;
output wire	F_BAR4;
output wire	F_BAR5;
output wire	F_BAR6;
output wire	F_BAR7;
output wire	USB_TX_BUSY_LED;
output wire	USB_RX_BUSY_LED;
output wire	5V_OUT_IDE_PORTS_RD-;
output wire	5V_OUT_IDE_PORTS_WR-;
output wire	VGA_R;
output wire	VGA_G;
output wire	VGA_B;
output wire	HSync;
output wire	VSync;
output wire	BUZZER;
output wire	F_BOARD_ACTIVE-;
output reg	FPGA_OUT_PRN_0;
output reg	FPGA_OUT_PRN_1;
output reg	FPGA_OUT_PRN_2;
output reg	FPGA_OUT_PRN_3;
output reg	FPGA_OUT_PRN_4;
output reg	FPGA_OUT_PRN_5;
output reg	FPGA_OUT_PRN_6;
output reg	FPGA_OUT_PRN_7;
output reg	FPGA_OUT_PRN_STROBE;
output wire	PRN_ACK_LED;
output wire	FPGA_OUT_PHANTOM;
output wire	S100_PHANTOM_LED;
output reg	RTC_CS;
output wire	RTC_SPI_SI;
output wire	RTC_SPI_CLK;
output wire	SD_CMD;
output wire	SD_CLK;
output wire	LED_4;
output wire	P1;
output wire	LED_1;
output wire	DIAG_LED;
output wire	SD_CS_B-;
output wire	FPGA_OUT_SPARE1;
output wire	SD_CS_A-;
output wire	FPGA_OUT_IDE_RD-;
output wire	FPGA_OUT_IDE_WR-;
output wire	FPGA_OUT_8255_SEL-;
output wire	FPGA_OUT_HIGH_ROM_LED-;
output wire	FPGA_OUT_LOW_ROM_LED-;
output wire	FPGA_OUT_HIGH_RAM_LED-;
output wire	LED_2;
output wire	LED_3;
inout wire	FPGA_BI_D0;
inout wire	FPGA_BI_D1;
inout wire	FPGA_BI_D2;
inout wire	FPGA_BI_D3;
inout wire	FPGA_BI_D4;
inout wire	FPGA_BI_D5;
inout wire	FPGA_BI_D6;
inout wire	FPGA_BI_D7;

wire	10mHz;
wire	25Mhz;
wire	2mHz;
wire	400_KHz_CLK;
wire	50mHz;
wire	ADDRESS_LATCH;
wire	BAR_IN_ENABLE-;
wire	BOARD_INT-;
wire	BOARD_WAIT-;
wire	[31:0] COUNTER_BUS;
wire	[31:0] CPU_CLK_COUNTER;
reg	[7:0] CTL;
wire	[7:0] CURSOR_X;
wire	[7:0] CURSOR_Y;
wire	[7:0] DATA_FROM_SDCARD;
wire	DATA_FROM_USB_PORT;
reg	DATA_IN_0_A;
reg	DATA_IN_1_A;
reg	DATA_IN_2_A;
reg	DATA_IN_3_A;
reg	DATA_IN_4_A;
reg	DATA_IN_5_A;
reg	DATA_IN_6_A;
reg	DATA_IN_7_A;
wire	DATA_OUT_D0;
wire	DATA_OUT_D1;
wire	DATA_OUT_D2;
wire	DATA_OUT_D3;
wire	DATA_OUT_D4;
wire	DATA_OUT_D5;
wire	DATA_OUT_D6;
wire	DATA_OUT_D7;
reg	[7:0] DATA_TO_SDCARD;
wire	DIP_5;
wire	DIP_6;
wire	DIP_7;
reg	DISABLE_ALL_ROM;
wire	END_SYNC;
wire	[11:0] FONT_A;
wire	[7:0] FONT_D;
wire	FORCE_LOW_SPEED-;
wire	FPGA_ROM;
wire	FPGA_ROM-;
wire	IDE_PORTA-;
wire	IDE_PORTB-;
wire	IDE_PORTC-;
wire	IDE_PORTCTRL-;
wire	IN_BOARD_RESET;
wire	IN_BOARD_RESET-;
wire	IN_CDSB-;
wire	IN_SDSB;
wire	IN_SDSB-;
wire	INTA_READ_DATA-;
wire	IO_INPUT;
wire	IO_OUTPUT;
wire	IOBYTE-;
wire	IOBYTE_OE-;
wire	JMP_ENABLE;
reg	JMP_ENABLE-;
wire	[15:0] LOCAL_ADDRESS_BUS;
wire	LOCAL_SD_SPI_CLK;
wire	MEM_READ;
wire	MEM_WRITE;
reg	[7:0] ocrx;
reg	[7:0] ocry;
wire	OUT_CPU_CLK;
wire	OUT_CPU_CLK-;
wire	OUT_MWRT;
wire	OUT_pDBIN;
wire	OUT_pWR-;
wire	OUT_RAM_READ-;
wire	OUT_RAM_WRITE-;
wire	OUT_sHLTA;
wire	OUT_sINP;
wire	OUT_sINTA;
wire	OUT_sM1;
wire	OUT_sMEMR;
wire	OUT_sOUT;
wire	OUT_sWO-;
wire	PORT_0-;
wire	PORT_1-;
wire	PORT_4-;
wire	PORT_5-;
wire	PORT_6-;
wire	PORT_7-;
wire	PORT_C0H-;
wire	PORT_C1H-;
wire	PORT_C2H-;
wire	PORT_C3H-;
wire	PORT_C4H-;
wire	PORT_C5H-;
wire	PORT_C6H-;
wire	PORT_C7H-;
wire	PORT_SELECT_68-;
wire	PORT_SELECT_69-;
wire	PORT_SELECT_6A-;
wire	PORT_SELECT_6B-;
wire	PORT_SELECT_6C-;
wire	PORT_SELECT_6D-;
wire	PORT_SELECT_6E-;
wire	PORT_SELECT_6F-;
wire	PRINTER_STATUS_PORT-;
wire	[6:0] PS2_ASCII_CODE;
wire	PS2_DATA-;
wire	PS2_DATA_IN;
reg	PS2_KEYBOARD_STATUS;
wire	PS2_STATUS-;
wire	PS2_STATUS_IN;
wire	pSYNC_RAW;
wire	[7:0] RAM_TEXT_D;
wire	READ_RAM;
reg	ROM_A12;
reg	ROM_A13;
wire	[13:0] ROM_ADDRESS;
wire	ROM_OE;
wire	S100_A0;
wire	S100_A1;
wire	S100_A10;
wire	S100_A11;
wire	S100_A12;
wire	S100_A13;
wire	S100_A14;
wire	S100_A15;
wire	S100_A16;
wire	S100_A17;
wire	S100_A18;
wire	S100_A19;
wire	S100_A2;
wire	S100_A3;
wire	S100_A4;
wire	S100_A5;
wire	S100_A6;
wire	S100_A7;
wire	S100_A8;
wire	S100_A9;
wire	S100_INT-;
wire	[31:0] SD_CARD_ADDRESS;
wire	SD_CARD_BUSY;
wire	[31:0] SD_CARD_CLK_DIV;
wire	SD_CARD_READ_DATA-;
reg	SD_READ;
wire	[1:0] SD_SLAVES;
reg	SD_WRITE;
reg	SDCARD_OUT_0;
reg	SDCARD_OUT_1;
reg	SDCARD_OUT_2;
reg	SDCARD_OUT_3;
reg	SDCARD_OUT_4;
reg	SDCARD_OUT_5;
reg	SDCARD_OUT_6;
reg	SDCARD_OUT_7;
wire	SERIAL_DATA_TO_USB_PORT;
wire	SPI_BUSY_FLAG;
wire	SPI_CLK;
wire	[31:0] SPI_CLK_DIV;
wire	[15:0] SPI_DATA_IN_BUS;
reg	[15:0] SPI_DATA_OUT_BUS;
wire	[31:0] SPI_INPUT_CS;
wire	SPI_MASTER_CLK;
reg	SPI_READ;
wire	SPI_RTC_READ_DATA-;
reg	SPI_SD_CLK_SPEED;
reg	SPI_WRITE;
reg	START_BUZZER;
wire	START_SYNC;
wire	STOP_BUZZER;
wire	[11:0] TEXT_A;
wire	UART_Busy;
wire	UART_Busy_Recieving;
wire	UART_Busy_Transmitting;
wire	UART_Byte_Recieved;
wire	UART_DATA_READY;
wire	UART_Error;
wire	USB_DATA-;
wire	USB_DATA_IN;
wire	USB_DATA_IN-;
wire	[7:0] USB_DATA_IN_BUS;
wire	USB_DATA_OUT;
reg	[7:0] USB_DATA_OUT_BUS;
wire	USB_STATUS-;
wire	USB_STATUS_IN;
wire	USB_STATUS_IN-;
wire	VGA_CURSOR_OE-;
wire	VGA_RAM_READ_DATA;
wire	VGA_RAM_READ_DATA-;
wire	VGA_RAM_SELECT;
wire	VGA_RAM_WRITE_DATA;
wire	WRITE;
wire	WRITE_RAM;
wire	[15:0] Z80_ADDRESS;
wire	Z80_BUSAK-;
reg	Z80_BUSRQ-;
wire	Z80_HALT-;
wire	Z80_INTA;
wire	Z80_IORQ;
wire	Z80_IORQ-;
wire	[7:0] Z80_LOCAL_D0;
wire	[7:0] Z80_LOCAL_DI;
wire	Z80_M1;
wire	Z80_M1-;
wire	Z80_MREQ;
wire	Z80_MREQ-;
wire	Z80_RD;
wire	Z80_RD-;
wire	Z80_RFSH-;
wire	Z80_WR;
wire	Z80_WR-;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_622;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_623;
wire	SYNTHESIZED_WIRE_624;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_625;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
reg	DFF_inst102;
reg	SYNTHESIZED_WIRE_626;
wire	SYNTHESIZED_WIRE_627;
wire	SYNTHESIZED_WIRE_628;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_629;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_630;
wire	[0:7] SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_631;
wire	SYNTHESIZED_WIRE_632;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_633;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_634;
wire	SYNTHESIZED_WIRE_635;
wire	SYNTHESIZED_WIRE_84;
wire	[0:7] SYNTHESIZED_WIRE_85;
reg	[7:0] SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_636;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_637;
wire	SYNTHESIZED_WIRE_638;
wire	SYNTHESIZED_WIRE_100;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_105;
wire	[0:7] SYNTHESIZED_WIRE_106;
reg	SYNTHESIZED_WIRE_107;
reg	[6:0] SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_639;
wire	[0:4] SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_640;
wire	SYNTHESIZED_WIRE_641;
wire	SYNTHESIZED_WIRE_642;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_643;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_644;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_146;
wire	SYNTHESIZED_WIRE_149;
reg	SYNTHESIZED_WIRE_154;
reg	SYNTHESIZED_WIRE_645;
wire	[7:0] SYNTHESIZED_WIRE_156;
reg	SYNTHESIZED_WIRE_646;
reg	SYNTHESIZED_WIRE_647;
reg	SYNTHESIZED_WIRE_648;
wire	SYNTHESIZED_WIRE_160;
wire	SYNTHESIZED_WIRE_649;
wire	SYNTHESIZED_WIRE_163;
reg	SYNTHESIZED_WIRE_650;
reg	SYNTHESIZED_WIRE_651;
reg	SYNTHESIZED_WIRE_652;
reg	SYNTHESIZED_WIRE_653;
wire	SYNTHESIZED_WIRE_168;
wire	SYNTHESIZED_WIRE_169;
wire	SYNTHESIZED_WIRE_654;
wire	SYNTHESIZED_WIRE_171;
wire	SYNTHESIZED_WIRE_173;
wire	SYNTHESIZED_WIRE_655;
wire	SYNTHESIZED_WIRE_656;
wire	SYNTHESIZED_WIRE_657;
wire	SYNTHESIZED_WIRE_658;
wire	SYNTHESIZED_WIRE_659;
wire	SYNTHESIZED_WIRE_660;
wire	SYNTHESIZED_WIRE_661;
wire	[0:1] SYNTHESIZED_WIRE_662;
wire	SYNTHESIZED_WIRE_199;
wire	[0:7] SYNTHESIZED_WIRE_200;
wire	SYNTHESIZED_WIRE_201;
wire	SYNTHESIZED_WIRE_663;
wire	SYNTHESIZED_WIRE_217;
wire	[0:7] SYNTHESIZED_WIRE_218;
reg	SYNTHESIZED_WIRE_219;
reg	SYNTHESIZED_WIRE_220;
reg	SYNTHESIZED_WIRE_221;
reg	SYNTHESIZED_WIRE_222;
reg	SYNTHESIZED_WIRE_223;
reg	SYNTHESIZED_WIRE_224;
reg	SYNTHESIZED_WIRE_225;
reg	SYNTHESIZED_WIRE_226;
wire	SYNTHESIZED_WIRE_227;
wire	SYNTHESIZED_WIRE_228;
wire	[0:7] SYNTHESIZED_WIRE_664;
wire	SYNTHESIZED_WIRE_665;
wire	SYNTHESIZED_WIRE_666;
wire	SYNTHESIZED_WIRE_667;
wire	SYNTHESIZED_WIRE_238;
wire	SYNTHESIZED_WIRE_239;
reg	SYNTHESIZED_WIRE_668;
wire	SYNTHESIZED_WIRE_240;
wire	[7:0] SYNTHESIZED_WIRE_242;
wire	SYNTHESIZED_WIRE_243;
wire	SYNTHESIZED_WIRE_244;
wire	SYNTHESIZED_WIRE_245;
wire	SYNTHESIZED_WIRE_246;
wire	[0:6] SYNTHESIZED_WIRE_669;
wire	SYNTHESIZED_WIRE_254;
wire	SYNTHESIZED_WIRE_255;
wire	SYNTHESIZED_WIRE_256;
wire	SYNTHESIZED_WIRE_257;
wire	SYNTHESIZED_WIRE_670;
wire	SYNTHESIZED_WIRE_259;
wire	SYNTHESIZED_WIRE_671;
wire	SYNTHESIZED_WIRE_262;
wire	SYNTHESIZED_WIRE_263;
wire	SYNTHESIZED_WIRE_264;
wire	SYNTHESIZED_WIRE_265;
wire	SYNTHESIZED_WIRE_672;
wire	SYNTHESIZED_WIRE_269;
wire	SYNTHESIZED_WIRE_270;
wire	SYNTHESIZED_WIRE_673;
wire	SYNTHESIZED_WIRE_674;
wire	SYNTHESIZED_WIRE_283;
wire	SYNTHESIZED_WIRE_284;
wire	[0:2] SYNTHESIZED_WIRE_285;
wire	SYNTHESIZED_WIRE_286;
wire	SYNTHESIZED_WIRE_675;
wire	SYNTHESIZED_WIRE_676;
wire	SYNTHESIZED_WIRE_293;
wire	SYNTHESIZED_WIRE_294;
wire	SYNTHESIZED_WIRE_677;
wire	SYNTHESIZED_WIRE_297;
wire	SYNTHESIZED_WIRE_678;
reg	DFF_inst143;
wire	SYNTHESIZED_WIRE_305;
wire	SYNTHESIZED_WIRE_306;
wire	SYNTHESIZED_WIRE_307;
wire	SYNTHESIZED_WIRE_309;
wire	SYNTHESIZED_WIRE_311;
reg	DFF_inst336;
wire	SYNTHESIZED_WIRE_679;
wire	SYNTHESIZED_WIRE_313;
wire	SYNTHESIZED_WIRE_680;
reg	SYNTHESIZED_WIRE_681;
wire	SYNTHESIZED_WIRE_316;
wire	SYNTHESIZED_WIRE_682;
wire	SYNTHESIZED_WIRE_319;
wire	SYNTHESIZED_WIRE_320;
wire	SYNTHESIZED_WIRE_322;
wire	SYNTHESIZED_WIRE_323;
wire	SYNTHESIZED_WIRE_324;
wire	SYNTHESIZED_WIRE_325;
reg	DFF_inst349;
wire	SYNTHESIZED_WIRE_327;
wire	SYNTHESIZED_WIRE_328;
reg	DFF_inst358;
wire	SYNTHESIZED_WIRE_330;
wire	SYNTHESIZED_WIRE_331;
wire	SYNTHESIZED_WIRE_332;
wire	SYNTHESIZED_WIRE_333;
wire	[0:31] SYNTHESIZED_WIRE_683;
wire	SYNTHESIZED_WIRE_336;
wire	SYNTHESIZED_WIRE_337;
wire	SYNTHESIZED_WIRE_338;
wire	SYNTHESIZED_WIRE_339;
wire	SYNTHESIZED_WIRE_340;
wire	SYNTHESIZED_WIRE_341;
wire	SYNTHESIZED_WIRE_342;
wire	SYNTHESIZED_WIRE_343;
wire	SYNTHESIZED_WIRE_344;
wire	SYNTHESIZED_WIRE_684;
wire	SYNTHESIZED_WIRE_685;
wire	SYNTHESIZED_WIRE_349;
wire	SYNTHESIZED_WIRE_686;
wire	SYNTHESIZED_WIRE_351;
wire	SYNTHESIZED_WIRE_687;
reg	DFF_inst377;
wire	SYNTHESIZED_WIRE_356;
wire	SYNTHESIZED_WIRE_357;
wire	SYNTHESIZED_WIRE_358;
wire	SYNTHESIZED_WIRE_688;
wire	SYNTHESIZED_WIRE_689;
wire	SYNTHESIZED_WIRE_690;
wire	SYNTHESIZED_WIRE_691;
wire	SYNTHESIZED_WIRE_372;
wire	SYNTHESIZED_WIRE_692;
reg	DFF_inst387;
wire	SYNTHESIZED_WIRE_377;
wire	SYNTHESIZED_WIRE_378;
wire	SYNTHESIZED_WIRE_379;
wire	SYNTHESIZED_WIRE_693;
wire	SYNTHESIZED_WIRE_381;
wire	SYNTHESIZED_WIRE_694;
wire	SYNTHESIZED_WIRE_695;
wire	SYNTHESIZED_WIRE_696;
wire	SYNTHESIZED_WIRE_697;
wire	SYNTHESIZED_WIRE_698;
wire	SYNTHESIZED_WIRE_699;
reg	SYNTHESIZED_WIRE_700;
wire	SYNTHESIZED_WIRE_701;
wire	SYNTHESIZED_WIRE_422;
wire	SYNTHESIZED_WIRE_426;
wire	SYNTHESIZED_WIRE_427;
wire	SYNTHESIZED_WIRE_702;
wire	SYNTHESIZED_WIRE_445;
wire	SYNTHESIZED_WIRE_703;
wire	SYNTHESIZED_WIRE_704;
wire	SYNTHESIZED_WIRE_462;
wire	SYNTHESIZED_WIRE_464;
wire	SYNTHESIZED_WIRE_465;
wire	SYNTHESIZED_WIRE_466;
wire	SYNTHESIZED_WIRE_467;
wire	SYNTHESIZED_WIRE_468;
wire	SYNTHESIZED_WIRE_469;
wire	SYNTHESIZED_WIRE_470;
wire	SYNTHESIZED_WIRE_705;
wire	SYNTHESIZED_WIRE_472;
wire	SYNTHESIZED_WIRE_476;
wire	SYNTHESIZED_WIRE_478;
wire	SYNTHESIZED_WIRE_479;
wire	SYNTHESIZED_WIRE_480;
wire	SYNTHESIZED_WIRE_481;
wire	SYNTHESIZED_WIRE_482;
wire	SYNTHESIZED_WIRE_483;
wire	SYNTHESIZED_WIRE_484;
wire	SYNTHESIZED_WIRE_706;
wire	SYNTHESIZED_WIRE_486;
wire	SYNTHESIZED_WIRE_707;
wire	SYNTHESIZED_WIRE_708;
wire	SYNTHESIZED_WIRE_709;
wire	SYNTHESIZED_WIRE_710;
wire	SYNTHESIZED_WIRE_711;
wire	SYNTHESIZED_WIRE_712;
reg	SYNTHESIZED_WIRE_497;
wire	SYNTHESIZED_WIRE_713;
reg	SYNTHESIZED_WIRE_500;
reg	SYNTHESIZED_WIRE_503;
wire	SYNTHESIZED_WIRE_505;
wire	SYNTHESIZED_WIRE_506;
reg	SYNTHESIZED_WIRE_714;
wire	SYNTHESIZED_WIRE_511;
wire	SYNTHESIZED_WIRE_715;
wire	SYNTHESIZED_WIRE_513;
wire	SYNTHESIZED_WIRE_716;
reg	SYNTHESIZED_WIRE_717;
wire	SYNTHESIZED_WIRE_535;
wire	SYNTHESIZED_WIRE_718;
wire	SYNTHESIZED_WIRE_719;
wire	SYNTHESIZED_WIRE_720;
reg	DFF_inst468;
wire	SYNTHESIZED_WIRE_559;
wire	SYNTHESIZED_WIRE_721;
wire	SYNTHESIZED_WIRE_722;
wire	SYNTHESIZED_WIRE_565;
wire	SYNTHESIZED_WIRE_723;
wire	SYNTHESIZED_WIRE_568;
wire	SYNTHESIZED_WIRE_569;
reg	DFF_inst512;
wire	[0:31] SYNTHESIZED_WIRE_724;
wire	SYNTHESIZED_WIRE_574;
wire	SYNTHESIZED_WIRE_575;
wire	SYNTHESIZED_WIRE_576;
wire	SYNTHESIZED_WIRE_577;
wire	SYNTHESIZED_WIRE_725;
wire	SYNTHESIZED_WIRE_581;
wire	SYNTHESIZED_WIRE_583;
wire	SYNTHESIZED_WIRE_586;
wire	SYNTHESIZED_WIRE_587;
wire	SYNTHESIZED_WIRE_588;
wire	SYNTHESIZED_WIRE_589;
wire	SYNTHESIZED_WIRE_590;
wire	SYNTHESIZED_WIRE_591;
wire	SYNTHESIZED_WIRE_726;
wire	SYNTHESIZED_WIRE_595;
reg	DFF_inst92;
wire	SYNTHESIZED_WIRE_727;
reg	DFF_inst97;
wire	SYNTHESIZED_WIRE_598;
wire	SYNTHESIZED_WIRE_599;
wire	SYNTHESIZED_WIRE_600;
wire	SYNTHESIZED_WIRE_603;
wire	[7:0] SYNTHESIZED_WIRE_604;
wire	SYNTHESIZED_WIRE_605;
wire	SYNTHESIZED_WIRE_606;
reg	DFF_inst95;
wire	SYNTHESIZED_WIRE_609;
wire	SYNTHESIZED_WIRE_728;
wire	SYNTHESIZED_WIRE_612;
wire	SYNTHESIZED_WIRE_613;
wire	SYNTHESIZED_WIRE_729;
wire	SYNTHESIZED_WIRE_615;
wire	SYNTHESIZED_WIRE_617;
wire	SYNTHESIZED_WIRE_730;

assign	FPGA_OUT_RAM_CS- = 0;
assign	FPGA_OUT_RAM_A17 = 0;
assign	FPGA_OUT_RAM_A18 = 0;
assign	LED_4 = SD_DO;
assign	FPGA_OUT_pHLDA = SYNTHESIZED_WIRE_625;
assign	PRN_ACK_LED = DFF_inst143;
assign	FPGA_OUT_PHANTOM = SYNTHESIZED_WIRE_283;
assign	P1 = SYNTHESIZED_WIRE_535;
assign	SD_CS_B- = SYNTHESIZED_WIRE_717;
assign	SD_CS_A- = SYNTHESIZED_WIRE_714;
assign	FPGA_OUT_IDE_RD- = SYNTHESIZED_WIRE_171;
assign	FPGA_OUT_IDE_WR- = SYNTHESIZED_WIRE_173;
assign	FPGA_OUT_8255_SEL- = SYNTHESIZED_WIRE_654;
assign	LED_2 = SYNTHESIZED_WIRE_714;
assign	LED_3 = SYNTHESIZED_WIRE_717;
assign	SYNTHESIZED_WIRE_1 = 1;
assign	SYNTHESIZED_WIRE_622 = 1;
assign	SYNTHESIZED_WIRE_623 = 0;
assign	SYNTHESIZED_WIRE_624 = 1;
assign	SYNTHESIZED_WIRE_19 = 1;
assign	SYNTHESIZED_WIRE_628 = 0;
assign	SYNTHESIZED_WIRE_629 = 1;
assign	SYNTHESIZED_WIRE_39 = 0;
assign	SYNTHESIZED_WIRE_44 = 1;
assign	SYNTHESIZED_WIRE_45 = 0;
assign	SYNTHESIZED_WIRE_55 = 0;
assign	SYNTHESIZED_WIRE_631 = 0;
assign	SYNTHESIZED_WIRE_632 = 1;
assign	SYNTHESIZED_WIRE_69 = 1;
assign	SYNTHESIZED_WIRE_634 = 0;
assign	SYNTHESIZED_WIRE_635 = 1;
assign	SYNTHESIZED_WIRE_85 = 1;
assign	SYNTHESIZED_WIRE_637 = 0;
assign	SYNTHESIZED_WIRE_106 = 1;
assign	SYNTHESIZED_WIRE_639 = 0;
assign	SYNTHESIZED_WIRE_120 = 0;
assign	SYNTHESIZED_WIRE_642 = 1;
assign	SYNTHESIZED_WIRE_644 = 1;
assign	SYNTHESIZED_WIRE_142 = 0;
assign	SYNTHESIZED_WIRE_144 = 0;
assign	SYNTHESIZED_WIRE_146 = 0;
assign	SYNTHESIZED_WIRE_657 = 1;
assign	SYNTHESIZED_WIRE_659 = 0;
assign	SYNTHESIZED_WIRE_660 = 1;
assign	SYNTHESIZED_WIRE_661 = 0;
assign	SYNTHESIZED_WIRE_662 = 0;
assign	SYNTHESIZED_WIRE_200 = 1;
assign	SYNTHESIZED_WIRE_218 = 1;
assign	SYNTHESIZED_WIRE_664 = 0;
assign	SYNTHESIZED_WIRE_239 = 1;
assign	SYNTHESIZED_WIRE_244 = 1;
assign	SYNTHESIZED_WIRE_246 = 1;
assign	SYNTHESIZED_WIRE_669 = 1;
assign	SYNTHESIZED_WIRE_671 = 1;
assign	SYNTHESIZED_WIRE_672 = 1;
assign	SYNTHESIZED_WIRE_673 = 0;
assign	SYNTHESIZED_WIRE_674 = 1;
assign	SYNTHESIZED_WIRE_285 = 1;
assign	SYNTHESIZED_WIRE_294 = 0;
assign	SYNTHESIZED_WIRE_678 = 1;
assign	SYNTHESIZED_WIRE_306 = 1;
assign	SYNTHESIZED_WIRE_307 = 0;
assign	SYNTHESIZED_WIRE_680 = 1;
assign	SYNTHESIZED_WIRE_682 = 1;
assign	SYNTHESIZED_WIRE_319 = 0;
assign	SYNTHESIZED_WIRE_322 = 1;
assign	SYNTHESIZED_WIRE_323 = 1;
assign	SYNTHESIZED_WIRE_327 = 1;
assign	SYNTHESIZED_WIRE_332 = 1;
assign	SYNTHESIZED_WIRE_683 = 1;
assign	SYNTHESIZED_WIRE_342 = 0;
assign	SYNTHESIZED_WIRE_684 = 1;
assign	SYNTHESIZED_WIRE_349 = 0;
assign	SYNTHESIZED_WIRE_687 = 1;
assign	SYNTHESIZED_WIRE_358 = 0;
assign	SYNTHESIZED_WIRE_689 = 0;
assign	SYNTHESIZED_WIRE_690 = 1;
assign	SYNTHESIZED_WIRE_692 = 1;
assign	SYNTHESIZED_WIRE_693 = 1;
assign	SYNTHESIZED_WIRE_695 = 1;
assign	SYNTHESIZED_WIRE_698 = 1;
assign	SYNTHESIZED_WIRE_699 = 0;
assign	SYNTHESIZED_WIRE_704 = 1;
assign	SYNTHESIZED_WIRE_705 = 0;
assign	SYNTHESIZED_WIRE_707 = 1;
assign	SYNTHESIZED_WIRE_711 = 1;
assign	SYNTHESIZED_WIRE_712 = 0;
assign	SYNTHESIZED_WIRE_715 = 1;
assign	SYNTHESIZED_WIRE_718 = 0;
assign	SYNTHESIZED_WIRE_723 = 1;
assign	SYNTHESIZED_WIRE_569 = 1;
assign	SYNTHESIZED_WIRE_724 = 1;
assign	SYNTHESIZED_WIRE_725 = 0;
assign	SYNTHESIZED_WIRE_609 = 1;
assign	SYNTHESIZED_WIRE_728 = 1;
assign	SYNTHESIZED_WIRE_612 = 1;
assign	SYNTHESIZED_WIRE_617 = 1;
assign	SYNTHESIZED_WIRE_730 = 1;




Microcomputer	b2v_inst(
	.n_reset(IN_BOARD_RESET-),
	.clk(OUT_CPU_CLK),
	.n_wait(SYNTHESIZED_WIRE_0),
	.n_int(BOARD_INT-),
	.n_nmi(SYNTHESIZED_WIRE_1),
	.n_busrq(Z80_BUSRQ-),
	.dataIn(Z80_LOCAL_DI),
	.n_wr(Z80_WR-),
	.n_rd(Z80_RD-),
	.n_mreq(Z80_MREQ-),
	.n_iorq(Z80_IORQ-),
	.n_busak(Z80_BUSAK-),
	.n_halt(Z80_HALT-),
	.n_rfsh(Z80_RFSH-),
	.n_m1(Z80_M1-),
	.address(Z80_ADDRESS),
	.dataOut(Z80_LOCAL_D0));


assign	pSYNC_RAW = ~(START_SYNC | END_SYNC | START_SYNC | SYNTHESIZED_WIRE_2);

assign	FPGA_ADD_OE- =  ~IN_SDSB-;

assign	FPGA_OUT_DO_OE- =  ~IN_SDSB-;


always@(posedge OUT_CPU_CLK or negedge SYNTHESIZED_WIRE_622 or negedge SYNTHESIZED_WIRE_622)
begin
if (!SYNTHESIZED_WIRE_622)
	begin
	DFF_inst102 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_622)
	begin
	DFF_inst102 <= 1;
	end
else
	begin
	DFF_inst102 <= SYNTHESIZED_WIRE_4;
	end
end


\74165 	b2v_inst103(
	.D(SYNTHESIZED_WIRE_623),
	.C(SYNTHESIZED_WIRE_624),
	.B(SYNTHESIZED_WIRE_624),
	.G(SYNTHESIZED_WIRE_623),
	.H(SYNTHESIZED_WIRE_623),
	.A(SYNTHESIZED_WIRE_624),
	.CLKIH(SYNTHESIZED_WIRE_623),
	.E(SYNTHESIZED_WIRE_623),
	.F(SYNTHESIZED_WIRE_623),
	.CLK(OUT_CPU_CLK-),
	.STLD(SYNTHESIZED_WIRE_15),
	.SER(SYNTHESIZED_WIRE_624),
	
	.QHN(SYNTHESIZED_WIRE_134));



assign	SYNTHESIZED_WIRE_2 =  ~Z80_RFSH-;

assign	FPGA_OUT_DI_OE- =  ~IN_SDSB-;


always@(posedge OUT_CPU_CLK- or negedge SYNTHESIZED_WIRE_625 or negedge SYNTHESIZED_WIRE_19)
begin
if (!SYNTHESIZED_WIRE_625)
	begin
	SYNTHESIZED_WIRE_626 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_19)
	begin
	SYNTHESIZED_WIRE_626 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_626 <= SYNTHESIZED_WIRE_625;
	end
end

assign	SYNTHESIZED_WIRE_4 = ~(SYNTHESIZED_WIRE_20 | FPGA_IN_pHOLD-);


assign	FPGA_OUT_CTL_DISABLE =  ~DFF_inst102;


assign	FPGA_OUT_STATUS_DISABLE =  ~SYNTHESIZED_WIRE_626;

assign	SYNTHESIZED_WIRE_625 =  ~Z80_BUSAK-;



\74373 	b2v_inst115(
	.D1(Z80_ADDRESS[0]),
	.D3(Z80_ADDRESS[2]),
	.D6(Z80_ADDRESS[5]),
	.D7(Z80_ADDRESS[6]),
	.D2(Z80_ADDRESS[1]),
	.G(ADDRESS_LATCH),
	.D4(Z80_ADDRESS[3]),
	.D5(Z80_ADDRESS[4]),
	.D8(Z80_ADDRESS[7]),
	.OEN(SYNTHESIZED_WIRE_627),
	.Q3(S100_A2),
	.Q6(S100_A5),
	.Q7(S100_A6),
	.Q2(S100_A1),
	.Q8(S100_A7),
	.Q4(S100_A3),
	.Q5(S100_A4),
	.Q1(S100_A0));


\74373 	b2v_inst116(
	.D1(Z80_ADDRESS[8]),
	.D3(Z80_ADDRESS[10]),
	.D6(Z80_ADDRESS[13]),
	.D7(Z80_ADDRESS[14]),
	.D2(Z80_ADDRESS[9]),
	.G(ADDRESS_LATCH),
	.D4(Z80_ADDRESS[11]),
	.D5(Z80_ADDRESS[12]),
	.D8(Z80_ADDRESS[15]),
	.OEN(SYNTHESIZED_WIRE_627),
	.Q3(SYNTHESIZED_WIRE_581),
	.Q6(SYNTHESIZED_WIRE_102),
	.Q7(SYNTHESIZED_WIRE_100),
	.Q2(SYNTHESIZED_WIRE_583),
	.Q8(SYNTHESIZED_WIRE_105),
	.Q4(SYNTHESIZED_WIRE_586),
	.Q5(SYNTHESIZED_WIRE_96),
	.Q1(SYNTHESIZED_WIRE_577));


\74373 	b2v_inst117(
	.D1(SYNTHESIZED_WIRE_628),
	.D3(SYNTHESIZED_WIRE_628),
	.D6(SYNTHESIZED_WIRE_628),
	.D7(SYNTHESIZED_WIRE_628),
	.D2(SYNTHESIZED_WIRE_628),
	.G(ADDRESS_LATCH),
	.D4(SYNTHESIZED_WIRE_628),
	.D5(SYNTHESIZED_WIRE_628),
	.D8(SYNTHESIZED_WIRE_628),
	.OEN(SYNTHESIZED_WIRE_627),
	.Q3(S100_A18),
	
	
	.Q2(S100_A17),
	
	.Q4(S100_A19),
	
	.Q1(S100_A16));

assign	SYNTHESIZED_WIRE_615 =  ~SYNTHESIZED_WIRE_32;



assign	SYNTHESIZED_WIRE_15 = ~(pSYNC_RAW & Z80_IORQ);


\74165 	b2v_inst121(
	.D(SYNTHESIZED_WIRE_629),
	.C(SYNTHESIZED_WIRE_629),
	.B(SYNTHESIZED_WIRE_629),
	.G(SYNTHESIZED_WIRE_629),
	.H(SYNTHESIZED_WIRE_629),
	.A(SYNTHESIZED_WIRE_629),
	.CLKIH(SYNTHESIZED_WIRE_39),
	.E(SYNTHESIZED_WIRE_629),
	.F(SYNTHESIZED_WIRE_629),
	.CLK(OUT_CPU_CLK-),
	.STLD(SYNTHESIZED_WIRE_42),
	.SER(SYNTHESIZED_WIRE_629),
	
	.QHN(SYNTHESIZED_WIRE_643));




always@(posedge IN_BOARD_RESET- or negedge SYNTHESIZED_WIRE_44 or negedge SYNTHESIZED_WIRE_46)
begin
if (!SYNTHESIZED_WIRE_44)
	begin
	JMP_ENABLE- <= 0;
	end
else
if (!SYNTHESIZED_WIRE_46)
	begin
	JMP_ENABLE- <= 1;
	end
else
	begin
	JMP_ENABLE- <= SYNTHESIZED_WIRE_45;
	end
end

assign	Z80_LOCAL_DI[0] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI0 : 1'bz;

assign	Z80_LOCAL_DI[1] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI1 : 1'bz;

assign	Z80_LOCAL_DI[2] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI2 : 1'bz;

assign	Z80_LOCAL_DI[3] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI3 : 1'bz;

assign	Z80_LOCAL_DI[4] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI4 : 1'bz;

assign	ADDRESS_LATCH = ~(pSYNC_RAW & OUT_CPU_CLK-);

assign	Z80_LOCAL_DI[5] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI5 : 1'bz;

assign	Z80_LOCAL_DI[6] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI6 : 1'bz;

assign	Z80_LOCAL_DI[7] = SYNTHESIZED_WIRE_630 ? FPGA_IN_DI7 : 1'bz;

assign	Z80_LOCAL_DI[7] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[0] : 1'bz;
assign	Z80_LOCAL_DI[6] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[1] : 1'bz;
assign	Z80_LOCAL_DI[5] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[2] : 1'bz;
assign	Z80_LOCAL_DI[4] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[3] : 1'bz;
assign	Z80_LOCAL_DI[3] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[4] : 1'bz;
assign	Z80_LOCAL_DI[2] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[5] : 1'bz;
assign	Z80_LOCAL_DI[1] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[6] : 1'bz;
assign	Z80_LOCAL_DI[0] = JMP_ENABLE ? SYNTHESIZED_WIRE_55[7] : 1'bz;

assign	FPGA_BI_D2 = WRITE_RAM ? DATA_OUT_D2 : 1'bz;

assign	Z80_LOCAL_DI[2] = READ_RAM ? FPGA_BI_D2 : 1'bz;

assign	FPGA_BI_D3 = WRITE_RAM ? DATA_OUT_D3 : 1'bz;

assign	Z80_LOCAL_DI[3] = READ_RAM ? FPGA_BI_D3 : 1'bz;


\74684 	b2v_inst138(
	.P2(SYNTHESIZED_WIRE_631),
	.Q2(SYNTHESIZED_WIRE_631),
	.P1(SYNTHESIZED_WIRE_631),
	.Q1(SYNTHESIZED_WIRE_631),
	.P0(SYNTHESIZED_WIRE_631),
	.Q0(SYNTHESIZED_WIRE_631),
	.P7(S100_A7),
	.Q7(SYNTHESIZED_WIRE_631),
	.Q6(SYNTHESIZED_WIRE_631),
	.P6(S100_A6),
	.Q5(SYNTHESIZED_WIRE_632),
	.P5(S100_A5),
	.P4(S100_A4),
	.Q4(SYNTHESIZED_WIRE_632),
	.Q3(SYNTHESIZED_WIRE_631),
	.P3(S100_A3),
	
	.EQUALN(SYNTHESIZED_WIRE_636));


assign	FPGA_OUT_HIGH_ROM_LED- = SYNTHESIZED_WIRE_67 | DISABLE_ALL_ROM;

assign	FPGA_BI_D4 = WRITE_RAM ? DATA_OUT_D4 : 1'bz;

assign	Z80_LOCAL_DI[4] = READ_RAM ? FPGA_BI_D4 : 1'bz;

assign	SYNTHESIZED_WIRE_667 = PORT_C1H- | SYNTHESIZED_WIRE_633;


always@(posedge IN_BOARD_RESET- or negedge FPGA_IN_PRN_ACK or negedge SYNTHESIZED_WIRE_70)
begin
if (!FPGA_IN_PRN_ACK)
	begin
	DFF_inst143 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_70)
	begin
	DFF_inst143 <= 1;
	end
else
	begin
	DFF_inst143 <= SYNTHESIZED_WIRE_69;
	end
end


assign	FPGA_BI_D5 = WRITE_RAM ? DATA_OUT_D5 : 1'bz;

assign	Z80_LOCAL_DI[5] = READ_RAM ? FPGA_BI_D5 : 1'bz;

assign	SYNTHESIZED_WIRE_238 = ~(IOBYTE- | SYNTHESIZED_WIRE_71);

assign	SYNTHESIZED_WIRE_283 = VGA_RAM_WRITE_DATA | VGA_RAM_READ_DATA;


\74684 	b2v_inst149(
	.P2(SYNTHESIZED_WIRE_634),
	.Q2(SYNTHESIZED_WIRE_634),
	.P1(SYNTHESIZED_WIRE_634),
	.Q1(SYNTHESIZED_WIRE_634),
	.P0(SYNTHESIZED_WIRE_634),
	.Q0(SYNTHESIZED_WIRE_634),
	.P7(S100_A15),
	.Q7(SYNTHESIZED_WIRE_635),
	.Q6(SYNTHESIZED_WIRE_635),
	.P6(S100_A14),
	.Q5(SYNTHESIZED_WIRE_635),
	.P5(S100_A13),
	.P4(S100_A12),
	.Q4(SYNTHESIZED_WIRE_635),
	.Q3(SYNTHESIZED_WIRE_634),
	.P3(SYNTHESIZED_WIRE_634),
	
	.EQUALN(SYNTHESIZED_WIRE_663));

assign	USB_TX_BUSY_LED =  ~UART_Busy;

assign	FPGA_BI_D6 = WRITE_RAM ? DATA_OUT_D6 : 1'bz;

assign	Z80_LOCAL_DI[6] = READ_RAM ? FPGA_BI_D6 : 1'bz;

assign	SYNTHESIZED_WIRE_84 =  ~UART_Busy_Transmitting;

assign	SYNTHESIZED_WIRE_331 = SYNTHESIZED_WIRE_84 & IN_BOARD_RESET-;


assign	FPGA_BI_D7 = WRITE_RAM ? DATA_OUT_D7 : 1'bz;

assign	Z80_LOCAL_DI[7] = READ_RAM ? FPGA_BI_D7 : 1'bz;



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_85 or USB_DATA_OUT or Z80_LOCAL_D0)
begin
if (~IN_BOARD_RESET-)
		USB_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_85)
		USB_DATA_OUT_BUS <= 1'b1;
else if (USB_DATA_OUT)
	USB_DATA_OUT_BUS <= Z80_LOCAL_D0;
end

assign	Z80_LOCAL_DI[7] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[7] : 1'bz;
assign	Z80_LOCAL_DI[6] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[6] : 1'bz;
assign	Z80_LOCAL_DI[5] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[5] : 1'bz;
assign	Z80_LOCAL_DI[4] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[4] : 1'bz;
assign	Z80_LOCAL_DI[3] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[3] : 1'bz;
assign	Z80_LOCAL_DI[2] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[2] : 1'bz;
assign	Z80_LOCAL_DI[1] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[1] : 1'bz;
assign	Z80_LOCAL_DI[0] = USB_DATA_IN ? SYNTHESIZED_WIRE_86[0] : 1'bz;


\74138 	b2v_inst16(
	.A(S100_A0),
	.B(S100_A1),
	.G1(SYNTHESIZED_WIRE_87),
	.C(S100_A2),
	.G2AN(SYNTHESIZED_WIRE_636),
	.G2BN(SYNTHESIZED_WIRE_636),
	.Y0N(IDE_PORTA-),
	.Y1N(IDE_PORTB-),
	.Y2N(IDE_PORTC-),
	.Y3N(IDE_PORTCTRL-),
	.Y4N(USB_STATUS-),
	.Y5N(USB_DATA-),
	.Y6N(IOBYTE-)
	);

assign	SYNTHESIZED_WIRE_264 = IN_BOARD_RESET- & PS2_DATA-;



ps2_keyboard_to_ascii	b2v_inst162(
	.clk(50mHz),
	.ps2_clk(FPGA_IN_PS2_CLK),
	.ps2_data(FPGA_IN_PS2_DATA),
	.ascii_new(SYNTHESIZED_WIRE_265),
	.ascii_code(PS2_ASCII_CODE));
	defparam	b2v_inst162.clk_freq = 50000000;
	defparam	b2v_inst162.ps2_debounce_counter_size = 8;

assign	SYNTHESIZED_WIRE_630 = SYNTHESIZED_WIRE_90 & SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_92 & IOBYTE_OE- & OUT_pDBIN & OUT_sINP & SYNTHESIZED_WIRE_93 & SYNTHESIZED_WIRE_94;

assign	USB_DATA_OUT = ~(USB_DATA- | OUT_pWR-);

assign	SYNTHESIZED_WIRE_305 = ~(SYNTHESIZED_WIRE_95 | OUT_pWR- | PORT_7-);

assign	SYNTHESIZED_WIRE_655 = FPGA_IN_PRN_ACK & IN_BOARD_RESET-;

assign	SYNTHESIZED_WIRE_257 = DIP_7 & FORCE_LOW_SPEED-;


\74157 	b2v_inst168(
	.A1(SYNTHESIZED_WIRE_96),
	.B1(SYNTHESIZED_WIRE_637),
	.SEL(SYNTHESIZED_WIRE_638),
	.B2(SYNTHESIZED_WIRE_637),
	.A3(SYNTHESIZED_WIRE_100),
	.B3(SYNTHESIZED_WIRE_637),
	.A2(SYNTHESIZED_WIRE_102),
	.B4(SYNTHESIZED_WIRE_637),
	.GN(SYNTHESIZED_WIRE_637),
	.A4(SYNTHESIZED_WIRE_105),
	.Y2(S100_A13),
	.Y1(S100_A12),
	.Y4(S100_A15),
	.Y3(S100_A14));


assign	SYNTHESIZED_WIRE_640 =  ~OUT_pDBIN;


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_106 or USB_DATA_IN or USB_DATA_IN_BUS)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_86 <= 1'b0;
else if (~SYNTHESIZED_WIRE_106)
		SYNTHESIZED_WIRE_86 <= 1'b1;
else if (USB_DATA_IN)
	SYNTHESIZED_WIRE_86 <= USB_DATA_IN_BUS;
end


assign	Z80_LOCAL_DI[0] = PS2_STATUS_IN ? SYNTHESIZED_WIRE_107 : 1'bz;

assign	Z80_LOCAL_DI[6] = PS2_DATA_IN ? SYNTHESIZED_WIRE_108[6] : 1'bz;
assign	Z80_LOCAL_DI[5] = PS2_DATA_IN ? SYNTHESIZED_WIRE_108[5] : 1'bz;
assign	Z80_LOCAL_DI[4] = PS2_DATA_IN ? SYNTHESIZED_WIRE_108[4] : 1'bz;
assign	Z80_LOCAL_DI[3] = PS2_DATA_IN ? SYNTHESIZED_WIRE_108[3] : 1'bz;
assign	Z80_LOCAL_DI[2] = PS2_DATA_IN ? SYNTHESIZED_WIRE_108[2] : 1'bz;
assign	Z80_LOCAL_DI[1] = PS2_DATA_IN ? SYNTHESIZED_WIRE_108[1] : 1'bz;
assign	Z80_LOCAL_DI[0] = PS2_DATA_IN ? SYNTHESIZED_WIRE_108[0] : 1'bz;


assign	SYNTHESIZED_WIRE_160 = OUT_sINP | OUT_sOUT;


\74684 	b2v_inst176(
	.P2(SYNTHESIZED_WIRE_639),
	.Q2(SYNTHESIZED_WIRE_639),
	.P1(SYNTHESIZED_WIRE_639),
	.Q1(SYNTHESIZED_WIRE_639),
	.P0(SYNTHESIZED_WIRE_639),
	.Q0(SYNTHESIZED_WIRE_639),
	.P7(S100_A7),
	.Q7(SYNTHESIZED_WIRE_639),
	.Q6(SYNTHESIZED_WIRE_639),
	.P6(S100_A6),
	.Q5(SYNTHESIZED_WIRE_639),
	.P5(S100_A5),
	.P4(S100_A4),
	.Q4(SYNTHESIZED_WIRE_639),
	.Q3(SYNTHESIZED_WIRE_639),
	.P3(S100_A3),
	
	.EQUALN(SYNTHESIZED_WIRE_649));

assign	SYNTHESIZED_WIRE_627 =  ~IN_SDSB-;

assign	SYNTHESIZED_WIRE_591 =  ~IN_SDSB-;

assign	CTL[7:3] =  ~SYNTHESIZED_WIRE_120;


\74373 	b2v_inst18(
	.D1(DIP7),
	.D3(DIP5),
	.D6(DIP_5),
	.D7(DIP_6),
	.D2(DIP6),
	.G(SYNTHESIZED_WIRE_640),
	.D4(DIP4),
	.D5(DIP3),
	.D8(DIP_7),
	.OEN(IOBYTE_OE-),
	.Q3(Z80_LOCAL_DI[2]),
	.Q6(Z80_LOCAL_DI[5]),
	.Q7(Z80_LOCAL_DI[6]),
	.Q2(Z80_LOCAL_DI[1]),
	.Q8(Z80_LOCAL_DI[7]),
	.Q4(Z80_LOCAL_DI[3]),
	.Q5(Z80_LOCAL_DI[4]),
	.Q1(Z80_LOCAL_DI[0]));




always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[0])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_645 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_645 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_645 <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[1])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_646 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_646 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_646 <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[2])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_647 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_647 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_647 <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[3])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_648 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_648 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_648 <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[4])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_650 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_650 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_650 <= Z80_LOCAL_D0;
end

assign	SYNTHESIZED_WIRE_163 =  ~OUT_sOUT;


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[5])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_652 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_652 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_652 <= Z80_LOCAL_D0;
end

assign	SYNTHESIZED_WIRE_137 =  ~OUT_pDBIN;

assign	BOARD_WAIT- = ~(SYNTHESIZED_WIRE_134 | SYNTHESIZED_WIRE_643 | SYNTHESIZED_WIRE_643);

assign	USB_DATA_IN = ~(USB_DATA- | SYNTHESIZED_WIRE_137);

assign	SYNTHESIZED_WIRE_149 =  ~OUT_pDBIN;


assign	UART_Busy = UART_Busy_Transmitting | UART_Busy_Transmitting;


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or UART_DATA_READY)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_221 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_221 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_221 <= UART_DATA_READY;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or UART_Busy)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_219 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_219 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_219 <= UART_Busy;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or UART_Byte_Recieved)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_222 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_222 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_222 <= UART_Byte_Recieved;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or UART_Busy_Recieving)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_220 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_220 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_220 <= UART_Busy_Recieving;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or SYNTHESIZED_WIRE_142)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_224 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_224 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_224 <= SYNTHESIZED_WIRE_142;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or SYNTHESIZED_WIRE_144)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_226 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_226 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_226 <= SYNTHESIZED_WIRE_144;
end

assign	WRITE_RAM = ~(JMP_ENABLE | OUT_RAM_WRITE-);



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or SYNTHESIZED_WIRE_146)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_223 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_223 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_223 <= SYNTHESIZED_WIRE_146;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_644 or USB_STATUS_IN or UART_Error)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_225 <= 1'b0;
else if (~SYNTHESIZED_WIRE_644)
		SYNTHESIZED_WIRE_225 <= 1'b1;
else if (USB_STATUS_IN)
	SYNTHESIZED_WIRE_225 <= UART_Error;
end



assign	SYNTHESIZED_WIRE_87 = OUT_sINP | OUT_sOUT;

assign	USB_STATUS_IN = ~(USB_STATUS- | SYNTHESIZED_WIRE_149);

assign	USB_STATUS_IN- =  ~USB_STATUS_IN;

assign	SYNTHESIZED_WIRE_513 = OUT_sINP | OUT_sOUT;


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[6])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_651 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_651 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_651 <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_642 or SYNTHESIZED_WIRE_641 or Z80_LOCAL_D0[7])
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_653 <= 1'b0;
else if (~SYNTHESIZED_WIRE_642)
		SYNTHESIZED_WIRE_653 <= 1'b1;
else if (SYNTHESIZED_WIRE_641)
	SYNTHESIZED_WIRE_653 <= Z80_LOCAL_D0;
end


assign	Z80_LOCAL_DI[7] = PS2_DATA_IN ? SYNTHESIZED_WIRE_154 : 1'bz;


assign	F_BAR0 =  ~SYNTHESIZED_WIRE_645;

assign	Z80_LOCAL_DI[7] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[7] : 1'bz;
assign	Z80_LOCAL_DI[6] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[6] : 1'bz;
assign	Z80_LOCAL_DI[5] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[5] : 1'bz;
assign	Z80_LOCAL_DI[4] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[4] : 1'bz;
assign	Z80_LOCAL_DI[3] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[3] : 1'bz;
assign	Z80_LOCAL_DI[2] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[2] : 1'bz;
assign	Z80_LOCAL_DI[1] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[1] : 1'bz;
assign	Z80_LOCAL_DI[0] = VGA_RAM_READ_DATA ? SYNTHESIZED_WIRE_156[0] : 1'bz;

assign	F_BAR1 =  ~SYNTHESIZED_WIRE_646;

assign	F_BAR2 =  ~SYNTHESIZED_WIRE_647;

assign	F_BAR3 =  ~SYNTHESIZED_WIRE_648;


\74138 	b2v_inst217(
	.A(S100_A0),
	.B(S100_A1),
	.G1(SYNTHESIZED_WIRE_160),
	.C(S100_A2),
	.G2AN(SYNTHESIZED_WIRE_649),
	.G2BN(SYNTHESIZED_WIRE_649),
	.Y0N(PORT_0-),
	
	.Y2N(PS2_STATUS-),
	.Y3N(PS2_DATA-),
	
	
	.Y6N(PORT_6-),
	.Y7N(PORT_7-));

assign	SYNTHESIZED_WIRE_641 = ~(OUT_pWR- | SYNTHESIZED_WIRE_163 | PORT_6-);

assign	F_BAR4 =  ~SYNTHESIZED_WIRE_650;

assign	USB_RX_BUSY_LED =  ~UART_Byte_Recieved;

assign	F_BAR6 =  ~SYNTHESIZED_WIRE_651;

assign	F_BAR5 =  ~SYNTHESIZED_WIRE_652;

assign	F_BAR7 =  ~SYNTHESIZED_WIRE_653;

assign	SYNTHESIZED_WIRE_46 = ~(MEM_READ & SYNTHESIZED_WIRE_168);

assign	SYNTHESIZED_WIRE_173 = ~(SYNTHESIZED_WIRE_169 & OUT_sOUT);

assign	SYNTHESIZED_WIRE_171 = ~(OUT_sINP & OUT_pDBIN);

assign	SYNTHESIZED_WIRE_169 =  ~OUT_pWR-;

assign	SYNTHESIZED_WIRE_654 = IDE_PORTA- & IDE_PORTB- & IDE_PORTC- & IDE_PORTCTRL-;

assign	5V_OUT_IDE_PORTS_RD- = SYNTHESIZED_WIRE_654 | SYNTHESIZED_WIRE_171;

assign	5V_OUT_IDE_PORTS_WR- = SYNTHESIZED_WIRE_654 | SYNTHESIZED_WIRE_173;

assign	DATA_OUT_D0 = Z80_LOCAL_D0[0] | Z80_LOCAL_D0[0];



always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[0])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_0 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_0 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_0 <= Z80_LOCAL_D0;
end

assign	SYNTHESIZED_WIRE_676 = PORT_C2H- | SYNTHESIZED_WIRE_658;


always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[1])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_1 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_1 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_1 <= Z80_LOCAL_D0;
end


always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[2])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_2 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_2 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_2 <= Z80_LOCAL_D0;
end


\74684 	b2v_inst235(
	.P2(SYNTHESIZED_WIRE_659),
	.Q2(SYNTHESIZED_WIRE_659),
	.P1(SYNTHESIZED_WIRE_659),
	.Q1(SYNTHESIZED_WIRE_659),
	.P0(SYNTHESIZED_WIRE_659),
	.Q0(SYNTHESIZED_WIRE_659),
	.P7(S100_A7),
	.Q7(SYNTHESIZED_WIRE_660),
	.Q6(SYNTHESIZED_WIRE_660),
	.P6(S100_A6),
	.Q5(SYNTHESIZED_WIRE_659),
	.P5(S100_A5),
	.P4(S100_A4),
	.Q4(SYNTHESIZED_WIRE_659),
	.Q3(SYNTHESIZED_WIRE_659),
	.P3(S100_A3),
	
	.EQUALN(SYNTHESIZED_WIRE_716));

assign	SYNTHESIZED_WIRE_633 =  ~OUT_pDBIN;

assign	CURSOR_X[7] = SYNTHESIZED_WIRE_661 | SYNTHESIZED_WIRE_661;

assign	CURSOR_Y[7:6] = SYNTHESIZED_WIRE_662 | SYNTHESIZED_WIRE_662;


assign	DATA_OUT_D1 = Z80_LOCAL_D0[1] | Z80_LOCAL_D0[1];


FPGA_ROM	b2v_inst240(
	.clock(25Mhz),
	.address(FONT_A),
	.q(FONT_D));

assign	IN_BOARD_RESET =  ~IN_BOARD_RESET-;



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_200 or SYNTHESIZED_WIRE_199 or Z80_LOCAL_D0)
begin
if (~IN_BOARD_RESET-)
		ocrx <= 1'b0;
else if (~SYNTHESIZED_WIRE_200)
		ocrx <= 1'b1;
else if (SYNTHESIZED_WIRE_199)
	ocrx <= Z80_LOCAL_D0;
end


assign	SYNTHESIZED_WIRE_201 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_199 = ~(OUT_pWR- | SYNTHESIZED_WIRE_201 | PORT_C0H-);


assign	SYNTHESIZED_WIRE_168 =  ~SYNTHESIZED_WIRE_663;


always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[3])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_3 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_3 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_3 <= Z80_LOCAL_D0;
end

assign	DATA_OUT_D2 = Z80_LOCAL_D0[2] | Z80_LOCAL_D0[2];


Counter01_32	b2v_inst250(
	.clock(OUT_CPU_CLK),
	.q(CPU_CLK_COUNTER));


always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[4])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_4 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_4 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_4 <= Z80_LOCAL_D0;
end


\74244 	b2v_inst252(
	.1A2(SYNTHESIZED_WIRE_646),
	.1A4(SYNTHESIZED_WIRE_648),
	.1A1(SYNTHESIZED_WIRE_645),
	.1A3(SYNTHESIZED_WIRE_647),
	.1GN(BAR_IN_ENABLE-),
	.2A3(SYNTHESIZED_WIRE_651),
	.2GN(BAR_IN_ENABLE-),
	.2A1(SYNTHESIZED_WIRE_650),
	.2A4(SYNTHESIZED_WIRE_653),
	.2A2(SYNTHESIZED_WIRE_652),
	.1Y2(Z80_LOCAL_DI[1]),
	.1Y4(Z80_LOCAL_DI[3]),
	.2Y1(Z80_LOCAL_DI[4]),
	.1Y1(Z80_LOCAL_DI[0]),
	.2Y3(Z80_LOCAL_DI[6]),
	.2Y4(Z80_LOCAL_DI[7]),
	.1Y3(Z80_LOCAL_DI[2]),
	.2Y2(Z80_LOCAL_DI[5]));


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_218 or SYNTHESIZED_WIRE_217 or Z80_LOCAL_D0)
begin
if (~IN_BOARD_RESET-)
		ocry <= 1'b0;
else if (~SYNTHESIZED_WIRE_218)
		ocry <= 1'b1;
else if (SYNTHESIZED_WIRE_217)
	ocry <= Z80_LOCAL_D0;
end

assign	SYNTHESIZED_WIRE_227 =  ~PORT_6-;


\74244 	b2v_inst255(
	.1A2(SYNTHESIZED_WIRE_219),
	.1A4(SYNTHESIZED_WIRE_220),
	.1A1(SYNTHESIZED_WIRE_221),
	.1A3(SYNTHESIZED_WIRE_222),
	.1GN(USB_STATUS_IN-),
	.2A3(SYNTHESIZED_WIRE_223),
	.2GN(USB_STATUS_IN-),
	.2A1(SYNTHESIZED_WIRE_224),
	.2A4(SYNTHESIZED_WIRE_225),
	.2A2(SYNTHESIZED_WIRE_226),
	.1Y2(Z80_LOCAL_DI[1]),
	.1Y4(Z80_LOCAL_DI[3]),
	.2Y1(Z80_LOCAL_DI[4]),
	.1Y1(Z80_LOCAL_DI[0]),
	.2Y3(Z80_LOCAL_DI[6]),
	.2Y4(Z80_LOCAL_DI[7]),
	.1Y3(Z80_LOCAL_DI[2]),
	.2Y2(Z80_LOCAL_DI[5]));

assign	BAR_IN_ENABLE- = ~(OUT_pDBIN & OUT_sINP & SYNTHESIZED_WIRE_227);

assign	SYNTHESIZED_WIRE_228 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_217 = ~(OUT_pWR- | SYNTHESIZED_WIRE_228 | PORT_C1H-);

assign	SYNTHESIZED_WIRE_242 = SYNTHESIZED_WIRE_664 | SYNTHESIZED_WIRE_664;

assign	DATA_OUT_D3 = Z80_LOCAL_D0[3] | Z80_LOCAL_D0[3];


\74373b 	b2v_inst260(
	.G(SYNTHESIZED_WIRE_665),
	.OEN(SYNTHESIZED_WIRE_666),
	.D(CURSOR_X),
	.Q(Z80_LOCAL_DI));


\74373b 	b2v_inst261(
	.G(SYNTHESIZED_WIRE_633),
	.OEN(SYNTHESIZED_WIRE_667),
	.D(CURSOR_Y),
	.Q(Z80_LOCAL_DI));


always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[5])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_5 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_5 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_5 <= Z80_LOCAL_D0;
end


assign	SYNTHESIZED_WIRE_638 = OUT_sINP | OUT_sOUT;



always@(posedge SYNTHESIZED_WIRE_238 or negedge IN_BOARD_RESET- or negedge SYNTHESIZED_WIRE_239)
begin
if (!IN_BOARD_RESET-)
	begin
	SYNTHESIZED_WIRE_668 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_239)
	begin
	SYNTHESIZED_WIRE_668 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_668 <= Z80_LOCAL_D0[0];
	end
end

assign	SYNTHESIZED_WIRE_240 =  ~S100_A15;

assign	FPGA_OUT_RAM_A16 = SYNTHESIZED_WIRE_668 & SYNTHESIZED_WIRE_240;


assign	DATA_OUT_D4 = Z80_LOCAL_D0[4] | Z80_LOCAL_D0[4];

assign	FPGA_OUT_HIGH_RAM_LED- =  ~SYNTHESIZED_WIRE_668;


Two_Port_RAM	b2v_inst271(
	.wren_a(VGA_RAM_WRITE_DATA),
	.wren_b(SYNTHESIZED_WIRE_664),
	.clock_a(25Mhz),
	.clock_b(25Mhz),
	.address_a(LOCAL_ADDRESS_BUS[11:0]),
	.address_b(TEXT_A),
	.data_a(Z80_LOCAL_D0),
	.data_b(SYNTHESIZED_WIRE_242),
	.q_a(SYNTHESIZED_WIRE_156),
	.q_b(RAM_TEXT_D));


always@(posedge SYNTHESIZED_WIRE_243 or negedge IN_BOARD_RESET- or negedge SYNTHESIZED_WIRE_244)
begin
if (!IN_BOARD_RESET-)
	begin
	DISABLE_ALL_ROM <= 0;
	end
else
if (!SYNTHESIZED_WIRE_244)
	begin
	DISABLE_ALL_ROM <= 1;
	end
else
	begin
	DISABLE_ALL_ROM <= Z80_LOCAL_D0[1];
	end
end

assign	SYNTHESIZED_WIRE_445 =  ~OUT_sOUT;


always@(posedge SYNTHESIZED_WIRE_245 or negedge IN_BOARD_RESET- or negedge SYNTHESIZED_WIRE_246)
begin
if (!IN_BOARD_RESET-)
	begin
	ROM_A12 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_246)
	begin
	ROM_A12 <= 1;
	end
else
	begin
	ROM_A12 <= Z80_LOCAL_D0[0];
	end
end



always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[6])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_6 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_6 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_6 <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_669 or PS2_DATA_IN or PS2_ASCII_CODE)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_108 <= 1'b0;
else if (~SYNTHESIZED_WIRE_669)
		SYNTHESIZED_WIRE_108 <= 1'b1;
else if (PS2_DATA_IN)
	SYNTHESIZED_WIRE_108 <= PS2_ASCII_CODE;
end



always@(SYNTHESIZED_WIRE_655 or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_656 or Z80_LOCAL_D0[7])
begin
if (~SYNTHESIZED_WIRE_655)
		FPGA_OUT_PRN_7 <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_7 <= 1'b1;
else if (SYNTHESIZED_WIRE_656)
	FPGA_OUT_PRN_7 <= Z80_LOCAL_D0;
end

assign	DATA_OUT_D5 = Z80_LOCAL_D0[5] | Z80_LOCAL_D0[5];


\74373b 	b2v_inst280(
	.G(ADDRESS_LATCH),
	.OEN(SYNTHESIZED_WIRE_254),
	.D(Z80_ADDRESS[7:0]),
	.Q(LOCAL_ADDRESS_BUS[7:0]));

assign	SYNTHESIZED_WIRE_254 =  ~IN_SDSB-;


\74373b 	b2v_inst282(
	.G(ADDRESS_LATCH),
	.OEN(SYNTHESIZED_WIRE_255),
	.D(Z80_ADDRESS[15:8]),
	.Q(LOCAL_ADDRESS_BUS[15:8]));

assign	SYNTHESIZED_WIRE_255 =  ~IN_SDSB-;

assign	SYNTHESIZED_WIRE_259 = ~(OUT_MWRT & VGA_RAM_SELECT);

assign	SYNTHESIZED_WIRE_42 = ~(Z80_MREQ & SYNTHESIZED_WIRE_256 & pSYNC_RAW);

assign	SYNTHESIZED_WIRE_256 =  ~FPGA_ROM-;


\21mux 	b2v_inst287(
	.S(SYNTHESIZED_WIRE_257),
	.B(2mHz),
	.A(25Mhz),
	.Y(OUT_CPU_CLK));

assign	SYNTHESIZED_WIRE_427 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_71 =  ~IO_OUTPUT;

assign	SYNTHESIZED_WIRE_729 = ~(Z80_RD- & SYNTHESIZED_WIRE_670);

assign	VGA_RAM_WRITE_DATA = ~(SYNTHESIZED_WIRE_259 | OUT_pWR-);

assign	SYNTHESIZED_WIRE_20 =  ~SYNTHESIZED_WIRE_626;


always@(posedge OUT_CPU_CLK or negedge SYNTHESIZED_WIRE_671 or negedge SYNTHESIZED_WIRE_671)
begin
if (!SYNTHESIZED_WIRE_671)
	begin
	Z80_BUSRQ- <= 0;
	end
else
if (!SYNTHESIZED_WIRE_671)
	begin
	Z80_BUSRQ- <= 1;
	end
else
	begin
	Z80_BUSRQ- <= FPGA_IN_pHOLD-;
	end
end


assign	VGA_RAM_READ_DATA = ~(SYNTHESIZED_WIRE_262 | SYNTHESIZED_WIRE_263);


always@(posedge SYNTHESIZED_WIRE_265 or negedge SYNTHESIZED_WIRE_264 or negedge SYNTHESIZED_WIRE_672)
begin
if (!SYNTHESIZED_WIRE_264)
	begin
	PS2_KEYBOARD_STATUS <= 0;
	end
else
if (!SYNTHESIZED_WIRE_672)
	begin
	PS2_KEYBOARD_STATUS <= 1;
	end
else
	begin
	PS2_KEYBOARD_STATUS <= SYNTHESIZED_WIRE_672;
	end
end


assign	SYNTHESIZED_WIRE_309 =  ~OUT_sMEMR;

assign	SYNTHESIZED_WIRE_94 =  ~READ_RAM;

assign	SYNTHESIZED_WIRE_720 = FPGA_ROM- & SYNTHESIZED_WIRE_663 & Z80_MREQ & Z80_MREQ;

assign	SYNTHESIZED_WIRE_0 = FPGA_IN_XRDY & FPGA_IN_RDY & BOARD_WAIT-;

assign	Z80_WR =  ~Z80_WR-;

assign	SYNTHESIZED_WIRE_719 = ~(PORT_SELECT_6C- | OUT_pWR-);

assign	ROM_OE = SYNTHESIZED_WIRE_269 & OUT_pDBIN & FPGA_ROM;

assign	SYNTHESIZED_WIRE_262 = ~(OUT_sMEMR & VGA_RAM_SELECT);

assign	SYNTHESIZED_WIRE_263 =  ~OUT_pDBIN;


assign	ROM_ADDRESS[5] = S100_A5 | S100_A5;

assign	ROM_ADDRESS[4] = S100_A4 | S100_A4;

assign	ROM_ADDRESS[3] = S100_A3 | S100_A3;

assign	ROM_ADDRESS[2] = S100_A2 | S100_A2;

assign	ROM_ADDRESS[1] = S100_A1 | S100_A1;

assign	Z80_IORQ =  ~Z80_IORQ-;

assign	ROM_ADDRESS[0] = S100_A0 | S100_A0;

assign	ROM_ADDRESS[11] = S100_A11 | S100_A11;

assign	ROM_ADDRESS[10] = S100_A10 | S100_A10;

assign	ROM_ADDRESS[9] = S100_A9 | S100_A9;

assign	ROM_ADDRESS[8] = S100_A8 | S100_A8;

assign	ROM_ADDRESS[7] = S100_A7 | S100_A7;

assign	ROM_ADDRESS[6] = S100_A6 | S100_A6;

assign	ROM_ADDRESS[12] = ROM_A12 | ROM_A12;

assign	FPGA_ROM =  ~FPGA_ROM-;

assign	VGA_RAM_SELECT =  ~SYNTHESIZED_WIRE_270;

assign	Z80_RD =  ~Z80_RD-;



\74684 	b2v_inst321(
	.P2(SYNTHESIZED_WIRE_673),
	.Q2(SYNTHESIZED_WIRE_673),
	.P1(SYNTHESIZED_WIRE_673),
	.Q1(SYNTHESIZED_WIRE_673),
	.P0(SYNTHESIZED_WIRE_673),
	.Q0(SYNTHESIZED_WIRE_673),
	.P7(S100_A15),
	.Q7(SYNTHESIZED_WIRE_674),
	.Q6(SYNTHESIZED_WIRE_674),
	.P6(S100_A14),
	.Q5(SYNTHESIZED_WIRE_674),
	.P5(S100_A13),
	.P4(S100_A12),
	.Q4(SYNTHESIZED_WIRE_673),
	.Q3(SYNTHESIZED_WIRE_673),
	.P3(SYNTHESIZED_WIRE_673),
	
	.EQUALN(SYNTHESIZED_WIRE_270));

assign	S100_PHANTOM_LED =  ~SYNTHESIZED_WIRE_283;

assign	VGA_RAM_READ_DATA- =  ~VGA_RAM_READ_DATA;



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_285 or SYNTHESIZED_WIRE_284 or Z80_LOCAL_D0)
begin
if (~IN_BOARD_RESET-)
		CTL <= 1'b0;
else if (~SYNTHESIZED_WIRE_285)
		CTL <= 1'b1;
else if (SYNTHESIZED_WIRE_284)
	CTL <= Z80_LOCAL_D0;
end

assign	SYNTHESIZED_WIRE_286 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_269 =  ~pSYNC_RAW;

assign	SYNTHESIZED_WIRE_284 = ~(OUT_pWR- | SYNTHESIZED_WIRE_286 | PORT_C2H-);

assign	SYNTHESIZED_WIRE_67 =  ~SYNTHESIZED_WIRE_675;

assign	Z80_MREQ =  ~Z80_MREQ-;

assign	SYNTHESIZED_WIRE_658 =  ~OUT_pDBIN;


\74373b 	b2v_inst331(
	.G(SYNTHESIZED_WIRE_658),
	.OEN(SYNTHESIZED_WIRE_676),
	.D(CURSOR_Y),
	.Q(Z80_LOCAL_DI));

assign	VGA_CURSOR_OE- = SYNTHESIZED_WIRE_666 & SYNTHESIZED_WIRE_667 & SYNTHESIZED_WIRE_676;


\74138 	b2v_inst333(
	.A(S100_A0),
	.B(S100_A1),
	.G1(SYNTHESIZED_WIRE_293),
	.C(SYNTHESIZED_WIRE_294),
	.G2AN(SYNTHESIZED_WIRE_677),
	.G2BN(SYNTHESIZED_WIRE_677),
	.Y0N(PORT_SELECT_68-),
	.Y1N(PORT_SELECT_69-),
	.Y2N(PORT_SELECT_6A-),
	.Y3N(PORT_SELECT_6B-)
	
	
	
	);


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_657 or SYNTHESIZED_WIRE_297 or Z80_LOCAL_D0[0])
begin
if (~IN_BOARD_RESET-)
		FPGA_OUT_PRN_STROBE <= 1'b0;
else if (~SYNTHESIZED_WIRE_657)
		FPGA_OUT_PRN_STROBE <= 1'b1;
else if (SYNTHESIZED_WIRE_297)
	FPGA_OUT_PRN_STROBE <= Z80_LOCAL_D0;
end


\74244 	b2v_inst335(
	.1A2(FPGA_IN_PRN_BUSY),
	.1A4(SYNTHESIZED_WIRE_678),
	.1A1(DFF_inst143),
	.1A3(SYNTHESIZED_WIRE_678),
	.1GN(PRINTER_STATUS_PORT-),
	.2A3(SYNTHESIZED_WIRE_678),
	.2GN(PRINTER_STATUS_PORT-),
	.2A1(SYNTHESIZED_WIRE_678),
	.2A4(SYNTHESIZED_WIRE_678),
	.2A2(SYNTHESIZED_WIRE_678),
	.1Y2(Z80_LOCAL_DI[1]),
	.1Y4(Z80_LOCAL_DI[3]),
	.2Y1(Z80_LOCAL_DI[4]),
	.1Y1(Z80_LOCAL_DI[0]),
	.2Y3(Z80_LOCAL_DI[6]),
	.2Y4(Z80_LOCAL_DI[7]),
	.1Y3(Z80_LOCAL_DI[2]),
	.2Y2(Z80_LOCAL_DI[5]));


always@(posedge SYNTHESIZED_WIRE_305 or negedge IN_BOARD_RESET- or negedge SYNTHESIZED_WIRE_306)
begin
if (!IN_BOARD_RESET-)
	begin
	DFF_inst336 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_306)
	begin
	DFF_inst336 <= 1;
	end
else
	begin
	DFF_inst336 <= Z80_LOCAL_D0[7];
	end
end


assign	SYNTHESIZED_WIRE_95 =  ~OUT_sOUT;


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_669 or PS2_DATA_IN or SYNTHESIZED_WIRE_307)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_154 <= 1'b0;
else if (~SYNTHESIZED_WIRE_669)
		SYNTHESIZED_WIRE_154 <= 1'b1;
else if (PS2_DATA_IN)
	SYNTHESIZED_WIRE_154 <= SYNTHESIZED_WIRE_307;
end

assign	FPGA_ROM- = SYNTHESIZED_WIRE_309 | DISABLE_ALL_ROM | SYNTHESIZED_WIRE_663;

assign	SYNTHESIZED_WIRE_311 =  ~OUT_pDBIN;

assign	PS2_DATA_IN = ~(PS2_DATA- | SYNTHESIZED_WIRE_311);

assign	FORCE_LOW_SPEED- =  ~DFF_inst336;

assign	SYNTHESIZED_WIRE_316 = SPI_READ | SPI_WRITE;

assign	BUZZER =  ~START_BUZZER;


always@(posedge SYNTHESIZED_WIRE_313 or negedge SYNTHESIZED_WIRE_679 or negedge SYNTHESIZED_WIRE_680)
begin
if (!SYNTHESIZED_WIRE_679)
	begin
	START_BUZZER <= 0;
	end
else
if (!SYNTHESIZED_WIRE_680)
	begin
	START_BUZZER <= 1;
	end
else
	begin
	START_BUZZER <= SYNTHESIZED_WIRE_680;
	end
end

assign	F_BOARD_ACTIVE- = SYNTHESIZED_WIRE_681 & CPU_CLK_COUNTER[20];


spi_16bit_master	b2v_inst347(
	.clock(SPI_CLK),
	.reset_n(IN_BOARD_RESET-),
	.enable(SYNTHESIZED_WIRE_316),
	.cpol(SYNTHESIZED_WIRE_682),
	.cpha(SYNTHESIZED_WIRE_682),
	.cont(SYNTHESIZED_WIRE_319),
	.miso(RTC_SPI_SO),
	.addr(SPI_INPUT_CS),
	.clk_div(SPI_CLK_DIV),
	.tx_data(SPI_DATA_OUT_BUS),
	.sclk(SPI_MASTER_CLK),
	.mosi(RTC_SPI_SI),
	.busy(SPI_BUSY_FLAG),
	.rx_data(SPI_DATA_IN_BUS)
	);
	defparam	b2v_inst347.d_width = 16;
	defparam	b2v_inst347.slaves = 4;

assign	SYNTHESIZED_WIRE_656 = ~(OUT_pWR- | SYNTHESIZED_WIRE_320 | PORT_C7H-);


always@(posedge COUNTER_BUS[16] or negedge SYNTHESIZED_WIRE_679 or negedge SYNTHESIZED_WIRE_322)
begin
if (!SYNTHESIZED_WIRE_679)
	begin
	DFF_inst349 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_322)
	begin
	DFF_inst349 <= 1;
	end
else
	begin
	DFF_inst349 <= START_BUZZER;
	end
end

assign	SYNTHESIZED_WIRE_589 =  ~Z80_HALT-;



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_323 or PS2_STATUS_IN or PS2_KEYBOARD_STATUS)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_107 <= 1'b0;
else if (~SYNTHESIZED_WIRE_323)
		SYNTHESIZED_WIRE_107 <= 1'b1;
else if (PS2_STATUS_IN)
	SYNTHESIZED_WIRE_107 <= PS2_KEYBOARD_STATUS;
end

assign	SYNTHESIZED_WIRE_324 =  ~OUT_pDBIN;

assign	PS2_STATUS_IN = ~(PS2_STATUS- | SYNTHESIZED_WIRE_324);



assign	SYNTHESIZED_WIRE_320 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_297 = ~(OUT_pWR- | SYNTHESIZED_WIRE_325 | PORT_C6H-);


always@(posedge COUNTER_BUS[16] or negedge SYNTHESIZED_WIRE_679 or negedge SYNTHESIZED_WIRE_327)
begin
if (!SYNTHESIZED_WIRE_679)
	begin
	DFF_inst358 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_327)
	begin
	DFF_inst358 <= 1;
	end
else
	begin
	DFF_inst358 <= DFF_inst349;
	end
end

assign	PRINTER_STATUS_PORT- = ~(OUT_pDBIN & OUT_sINP & SYNTHESIZED_WIRE_328);

assign	Z80_M1 =  ~Z80_M1-;

assign	SYNTHESIZED_WIRE_328 =  ~PORT_C7H-;


assign	STOP_BUZZER =  ~DFF_inst358;

assign	SYNTHESIZED_WIRE_325 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_679 = IN_BOARD_RESET- & STOP_BUZZER;

assign	SYNTHESIZED_WIRE_70 =  ~SYNTHESIZED_WIRE_656;


assign	SYNTHESIZED_WIRE_313 = ~(OUT_pWR- | SYNTHESIZED_WIRE_330 | PORT_0-);

assign	SYNTHESIZED_WIRE_330 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_351 = ~(PORT_SELECT_6B- | OUT_pWR-);


\74164 	b2v_inst37(
	.CLRN(SYNTHESIZED_WIRE_331),
	.CLK(OUT_CPU_CLK),
	.B(SYNTHESIZED_WIRE_332),
	.A(USB_DATA_OUT),
	
	
	
	
	
	
	
	.QB(SYNTHESIZED_WIRE_606));

assign	SYNTHESIZED_WIRE_372 = ~(PORT_SELECT_6B- | SYNTHESIZED_WIRE_333);


assign	SPI_CLK_DIV =  ~SYNTHESIZED_WIRE_683;


assign	SPI_INPUT_CS =  ~SYNTHESIZED_WIRE_683;


\74148 	b2v_inst375(
	.5N(SYNTHESIZED_WIRE_336),
	.0N(SYNTHESIZED_WIRE_337),
	.1N(SYNTHESIZED_WIRE_338),
	.2N(SYNTHESIZED_WIRE_339),
	.3N(SYNTHESIZED_WIRE_340),
	.4N(SYNTHESIZED_WIRE_341),
	.EIN(SYNTHESIZED_WIRE_342),
	.6N(SYNTHESIZED_WIRE_343),
	.7N(SYNTHESIZED_WIRE_344),
	.A1N(SYNTHESIZED_WIRE_481),
	.A0N(SYNTHESIZED_WIRE_479),
	.A2N(SYNTHESIZED_WIRE_484),
	
	.GSN(SYNTHESIZED_WIRE_482));


\74373 	b2v_inst376(
	.D1(SYNTHESIZED_WIRE_684),
	.D3(RTC_INT),
	.D6(FPGA_IN_INT_B-),
	.D7(FPGA_IN_INT_A-),
	.D2(SYNTHESIZED_WIRE_684),
	.G(SYNTHESIZED_WIRE_685),
	.D4(FPGA_IN_INT_D-),
	.D5(FPGA_IN_INT_C-),
	.D8(SYNTHESIZED_WIRE_684),
	.OEN(SYNTHESIZED_WIRE_349),
	.Q3(SYNTHESIZED_WIRE_340),
	.Q6(SYNTHESIZED_WIRE_343),
	.Q7(SYNTHESIZED_WIRE_344),
	.Q2(SYNTHESIZED_WIRE_339),
	.Q8(SYNTHESIZED_WIRE_337),
	.Q4(SYNTHESIZED_WIRE_341),
	.Q5(SYNTHESIZED_WIRE_336),
	.Q1(SYNTHESIZED_WIRE_338));


always@(posedge SYNTHESIZED_WIRE_351 or negedge SYNTHESIZED_WIRE_686 or negedge SYNTHESIZED_WIRE_687)
begin
if (!SYNTHESIZED_WIRE_686)
	begin
	DFF_inst377 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_687)
	begin
	DFF_inst377 <= 1;
	end
else
	begin
	DFF_inst377 <= SYNTHESIZED_WIRE_687;
	end
end



always@(posedge SPI_CLK or negedge SYNTHESIZED_WIRE_686 or negedge SYNTHESIZED_WIRE_687)
begin
if (!SYNTHESIZED_WIRE_686)
	begin
	SPI_WRITE <= 0;
	end
else
if (!SYNTHESIZED_WIRE_687)
	begin
	SPI_WRITE <= 1;
	end
else
	begin
	SPI_WRITE <= DFF_inst377;
	end
end

assign	DATA_OUT_D6 = Z80_LOCAL_D0[6] | Z80_LOCAL_D0[6];

assign	SYNTHESIZED_WIRE_356 =  ~SPI_BUSY_FLAG;

assign	SYNTHESIZED_WIRE_686 = SYNTHESIZED_WIRE_356 & IN_BOARD_RESET-;

assign	SPI_CLK =  ~COUNTER_BUS[4];


assign	SYNTHESIZED_WIRE_333 =  ~OUT_pDBIN;


\74138 	b2v_inst385(
	.A(S100_A0),
	.B(S100_A1),
	.G1(SYNTHESIZED_WIRE_357),
	.C(SYNTHESIZED_WIRE_358),
	.G2AN(SYNTHESIZED_WIRE_688),
	.G2BN(SYNTHESIZED_WIRE_688),
	.Y0N(PORT_SELECT_6C-),
	.Y1N(PORT_SELECT_6D-),
	.Y2N(PORT_SELECT_6E-),
	.Y3N(PORT_SELECT_6F-)
	
	
	
	);


\74684 	b2v_inst386(
	.P2(S100_A2),
	.Q2(SYNTHESIZED_WIRE_689),
	.P1(SYNTHESIZED_WIRE_689),
	.Q1(SYNTHESIZED_WIRE_689),
	.P0(SYNTHESIZED_WIRE_689),
	.Q0(SYNTHESIZED_WIRE_689),
	.P7(S100_A7),
	.Q7(SYNTHESIZED_WIRE_689),
	.Q6(SYNTHESIZED_WIRE_690),
	.P6(S100_A6),
	.Q5(SYNTHESIZED_WIRE_690),
	.P5(S100_A5),
	.P4(S100_A4),
	.Q4(SYNTHESIZED_WIRE_689),
	.Q3(SYNTHESIZED_WIRE_690),
	.P3(S100_A3),
	
	.EQUALN(SYNTHESIZED_WIRE_677));


always@(posedge SYNTHESIZED_WIRE_372 or negedge SYNTHESIZED_WIRE_691 or negedge SYNTHESIZED_WIRE_692)
begin
if (!SYNTHESIZED_WIRE_691)
	begin
	DFF_inst387 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_692)
	begin
	DFF_inst387 <= 1;
	end
else
	begin
	DFF_inst387 <= SYNTHESIZED_WIRE_692;
	end
end



always@(posedge SPI_CLK or negedge SYNTHESIZED_WIRE_691 or negedge SYNTHESIZED_WIRE_692)
begin
if (!SYNTHESIZED_WIRE_691)
	begin
	SPI_READ <= 0;
	end
else
if (!SYNTHESIZED_WIRE_692)
	begin
	SPI_READ <= 1;
	end
else
	begin
	SPI_READ <= DFF_inst387;
	end
end

assign	DATA_OUT_D7 = Z80_LOCAL_D0[7] | Z80_LOCAL_D0[7];

assign	SYNTHESIZED_WIRE_377 =  ~SPI_BUSY_FLAG;

assign	SYNTHESIZED_WIRE_691 = SYNTHESIZED_WIRE_377 & IN_BOARD_RESET-;

assign	SYNTHESIZED_WIRE_702 = ~(OUT_pWR- | PORT_SELECT_68- | SYNTHESIZED_WIRE_378);



assign	SYNTHESIZED_WIRE_293 = OUT_sINP | OUT_sOUT;

assign	SYNTHESIZED_WIRE_378 =  ~OUT_sOUT;


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_379 or Z80_LOCAL_D0[0])
begin
if (~IN_BOARD_RESET-)
		RTC_CS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		RTC_CS <= 1'b1;
else if (SYNTHESIZED_WIRE_379)
	RTC_CS <= Z80_LOCAL_D0;
end

assign	SYNTHESIZED_WIRE_379 = ~(OUT_pWR- | PORT_SELECT_6A- | SYNTHESIZED_WIRE_381);

assign	SYNTHESIZED_WIRE_381 =  ~OUT_sOUT;


PLL01_50	b2v_inst4(
	.inclk0(50mHz),
	.c0(2mHz),
	.c1(400_KHz_CLK),
	.c2(10mHz),
	.c3(25Mhz));





always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[7])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_7_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_7_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_7_A <= SPI_DATA_IN_BUS;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[6])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_6_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_6_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_6_A <= SPI_DATA_IN_BUS;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[5])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_5_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_5_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_5_A <= SPI_DATA_IN_BUS;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[4])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_4_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_4_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_4_A <= SPI_DATA_IN_BUS;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[3])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_3_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_3_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_3_A <= SPI_DATA_IN_BUS;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[2])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_2_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_2_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_2_A <= SPI_DATA_IN_BUS;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[1])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_1_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_1_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_1_A <= SPI_DATA_IN_BUS;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_694 or SPI_DATA_IN_BUS[0])
begin
if (~IN_BOARD_RESET-)
		DATA_IN_0_A <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		DATA_IN_0_A <= 1'b1;
else if (SYNTHESIZED_WIRE_694)
	DATA_IN_0_A <= SPI_DATA_IN_BUS;
end

assign	READ_RAM =  ~OUT_RAM_READ-;


\74244 	b2v_inst410(
	.1A2(DATA_IN_6_A),
	.1A4(DATA_IN_4_A),
	.1A1(DATA_IN_7_A),
	.1A3(DATA_IN_5_A),
	.1GN(SYNTHESIZED_WIRE_696),
	.2A3(DATA_IN_1_A),
	.2GN(SYNTHESIZED_WIRE_696),
	.2A1(DATA_IN_3_A),
	.2A4(DATA_IN_0_A),
	.2A2(DATA_IN_2_A),
	.1Y2(Z80_LOCAL_DI[6]),
	.1Y4(Z80_LOCAL_DI[4]),
	.2Y1(Z80_LOCAL_DI[3]),
	.1Y1(Z80_LOCAL_DI[7]),
	.2Y3(Z80_LOCAL_DI[1]),
	.2Y4(Z80_LOCAL_DI[0]),
	.1Y3(Z80_LOCAL_DI[5]),
	.2Y2(Z80_LOCAL_DI[2]));


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_695 or SYNTHESIZED_WIRE_697 or SPI_BUSY_FLAG)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_700 <= 1'b0;
else if (~SYNTHESIZED_WIRE_695)
		SYNTHESIZED_WIRE_700 <= 1'b1;
else if (SYNTHESIZED_WIRE_697)
	SYNTHESIZED_WIRE_700 <= SPI_BUSY_FLAG;
end


\74684 	b2v_inst412(
	.P2(S100_A2),
	.Q2(SYNTHESIZED_WIRE_698),
	.P1(SYNTHESIZED_WIRE_699),
	.Q1(SYNTHESIZED_WIRE_699),
	.P0(SYNTHESIZED_WIRE_699),
	.Q0(SYNTHESIZED_WIRE_699),
	.P7(S100_A7),
	.Q7(SYNTHESIZED_WIRE_699),
	.Q6(SYNTHESIZED_WIRE_698),
	.P6(S100_A6),
	.Q5(SYNTHESIZED_WIRE_698),
	.P5(S100_A5),
	.P4(S100_A4),
	.Q4(SYNTHESIZED_WIRE_699),
	.Q3(SYNTHESIZED_WIRE_698),
	.P3(S100_A3),
	
	.EQUALN(SYNTHESIZED_WIRE_688));


\74244 	b2v_inst413(
	.1A2(SYNTHESIZED_WIRE_700),
	.1A4(SYNTHESIZED_WIRE_700),
	.1A1(SYNTHESIZED_WIRE_700),
	.1A3(SYNTHESIZED_WIRE_700),
	.1GN(SYNTHESIZED_WIRE_701),
	.2A3(SYNTHESIZED_WIRE_700),
	.2GN(SYNTHESIZED_WIRE_701),
	.2A1(SYNTHESIZED_WIRE_700),
	.2A4(SYNTHESIZED_WIRE_700),
	.2A2(SYNTHESIZED_WIRE_700),
	.1Y2(Z80_LOCAL_DI[6]),
	.1Y4(Z80_LOCAL_DI[4]),
	.2Y1(Z80_LOCAL_DI[3]),
	.1Y1(Z80_LOCAL_DI[7]),
	.2Y3(Z80_LOCAL_DI[1]),
	.2Y4(Z80_LOCAL_DI[0]),
	.1Y3(Z80_LOCAL_DI[5]),
	.2Y2(Z80_LOCAL_DI[2]));

assign	SYNTHESIZED_WIRE_694 = OUT_pDBIN & SYNTHESIZED_WIRE_422 & OUT_sINP;

assign	SYNTHESIZED_WIRE_422 =  ~PORT_SELECT_69-;

assign	SPI_RTC_READ_DATA- = ~(SYNTHESIZED_WIRE_694 | SYNTHESIZED_WIRE_697);

assign	SYNTHESIZED_WIRE_696 =  ~SYNTHESIZED_WIRE_694;

assign	SYNTHESIZED_WIRE_697 = OUT_pDBIN & SYNTHESIZED_WIRE_426 & OUT_sINP;

assign	SYNTHESIZED_WIRE_426 =  ~PORT_SELECT_6A-;

assign	SYNTHESIZED_WIRE_245 = ~(SYNTHESIZED_WIRE_427 | OUT_pWR- | PORT_7-);

assign	SYNTHESIZED_WIRE_701 =  ~SYNTHESIZED_WIRE_697;



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[7])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[6])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[5])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[4])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[3])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[2])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[1])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_693 or SYNTHESIZED_WIRE_702 or Z80_LOCAL_D0[0])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_693)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_702)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end

assign	SYNTHESIZED_WIRE_243 = ~(SYNTHESIZED_WIRE_445 | OUT_pWR- | PORT_7-);

assign	SYNTHESIZED_WIRE_92 = VGA_RAM_READ_DATA- & VGA_CURSOR_OE- & SPI_RTC_READ_DATA-;



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[7])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[6])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[5])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[4])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[3])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[2])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[1])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_704 or SYNTHESIZED_WIRE_703 or Z80_LOCAL_D0[0])
begin
if (~IN_BOARD_RESET-)
		SPI_DATA_OUT_BUS <= 1'b0;
else if (~SYNTHESIZED_WIRE_704)
		SPI_DATA_OUT_BUS <= 1'b1;
else if (SYNTHESIZED_WIRE_703)
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
end


FPGA_ROM_16K	b2v_inst44(
	.clock(ROM_OE),
	.address(ROM_ADDRESS),
	.q(SYNTHESIZED_WIRE_604));

assign	SYNTHESIZED_WIRE_703 = ~(OUT_pWR- | PORT_SELECT_69- | SYNTHESIZED_WIRE_462);

assign	SYNTHESIZED_WIRE_462 =  ~OUT_sOUT;



assign	SYNTHESIZED_WIRE_464 =  ~SYNTHESIZED_WIRE_685;

assign	SYNTHESIZED_WIRE_465 =  ~SYNTHESIZED_WIRE_464;

assign	SYNTHESIZED_WIRE_466 =  ~SYNTHESIZED_WIRE_465;

assign	SYNTHESIZED_WIRE_467 =  ~SYNTHESIZED_WIRE_466;

assign	SYNTHESIZED_WIRE_468 =  ~SYNTHESIZED_WIRE_467;

assign	SYNTHESIZED_WIRE_469 =  ~SYNTHESIZED_WIRE_468;

assign	FPGA_BI_D0 = WRITE_RAM ? DATA_OUT_D0 : 1'bz;

assign	SYNTHESIZED_WIRE_470 =  ~SYNTHESIZED_WIRE_469;

assign	SYNTHESIZED_WIRE_483 =  ~SYNTHESIZED_WIRE_470;


\74244 	b2v_inst452(
	.1A2(SYNTHESIZED_WIRE_705),
	.1A4(SYNTHESIZED_WIRE_472),
	.1A1(SYNTHESIZED_WIRE_705),
	.1A3(SYNTHESIZED_WIRE_705),
	.1GN(INTA_READ_DATA-),
	.2A3(SYNTHESIZED_WIRE_705),
	.2GN(INTA_READ_DATA-),
	.2A1(SYNTHESIZED_WIRE_476),
	.2A4(SYNTHESIZED_WIRE_705),
	.2A2(SYNTHESIZED_WIRE_478),
	.1Y2(Z80_LOCAL_DI[1]),
	.1Y4(Z80_LOCAL_DI[3]),
	.2Y1(Z80_LOCAL_DI[4]),
	.1Y1(Z80_LOCAL_DI[0]),
	.2Y3(Z80_LOCAL_DI[6]),
	.2Y4(Z80_LOCAL_DI[7]),
	.1Y3(Z80_LOCAL_DI[2]),
	.2Y2(Z80_LOCAL_DI[5]));

assign	SYNTHESIZED_WIRE_472 =  ~SYNTHESIZED_WIRE_479;

assign	SYNTHESIZED_WIRE_93 = PRINTER_STATUS_PORT- & INTA_READ_DATA-;

assign	BOARD_INT- = SYNTHESIZED_WIRE_480 & S100_INT-;

assign	SYNTHESIZED_WIRE_685 =  ~OUT_sINTA;

assign	SYNTHESIZED_WIRE_476 =  ~SYNTHESIZED_WIRE_481;

assign	SYNTHESIZED_WIRE_480 = FPGA_IN_ENABLE_INTA | SYNTHESIZED_WIRE_482;

assign	INTA_READ_DATA- = SYNTHESIZED_WIRE_483 | FPGA_IN_ENABLE_INTA;

assign	Z80_LOCAL_DI[0] = READ_RAM ? FPGA_BI_D0 : 1'bz;



assign	SYNTHESIZED_WIRE_478 =  ~SYNTHESIZED_WIRE_484;


assign	SYNTHESIZED_WIRE_357 = OUT_sINP | OUT_sOUT;

assign	SYNTHESIZED_WIRE_511 = ~(PORT_SELECT_6D- | OUT_pWR-);


assign	SYNTHESIZED_WIRE_721 = ~(PORT_SELECT_6E- | OUT_pWR-);


always@(posedge SYNTHESIZED_WIRE_486 or negedge SYNTHESIZED_WIRE_706 or negedge SYNTHESIZED_WIRE_707)
begin
if (!SYNTHESIZED_WIRE_706)
	begin
	DFF_inst468 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_707)
	begin
	DFF_inst468 <= 1;
	end
else
	begin
	DFF_inst468 <= SYNTHESIZED_WIRE_707;
	end
end


\74244 	b2v_inst469(
	.1A2(SDCARD_OUT_6),
	.1A4(SDCARD_OUT_4),
	.1A1(SDCARD_OUT_7),
	.1A3(SDCARD_OUT_5),
	.1GN(SYNTHESIZED_WIRE_708),
	.2A3(SDCARD_OUT_1),
	.2GN(SYNTHESIZED_WIRE_708),
	.2A1(SDCARD_OUT_3),
	.2A4(SDCARD_OUT_0),
	.2A2(SDCARD_OUT_2),
	.1Y2(Z80_LOCAL_DI[6]),
	.1Y4(Z80_LOCAL_DI[4]),
	.2Y1(Z80_LOCAL_DI[3]),
	.1Y1(Z80_LOCAL_DI[7]),
	.2Y3(Z80_LOCAL_DI[1]),
	.2Y4(Z80_LOCAL_DI[0]),
	.1Y3(Z80_LOCAL_DI[5]),
	.2Y2(Z80_LOCAL_DI[2]));

assign	FPGA_BI_D1 = WRITE_RAM ? DATA_OUT_D1 : 1'bz;

assign	SD_CARD_READ_DATA- = ~(SYNTHESIZED_WIRE_709 | SYNTHESIZED_WIRE_710);


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_710 or SD_CARD_BUSY)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_497 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SYNTHESIZED_WIRE_497 <= 1'b1;
else if (SYNTHESIZED_WIRE_710)
	SYNTHESIZED_WIRE_497 <= SD_CARD_BUSY;
end


\74244 	b2v_inst472(
	.1A2(SYNTHESIZED_WIRE_712),
	.1A4(SYNTHESIZED_WIRE_712),
	.1A1(SYNTHESIZED_WIRE_497),
	.1A3(SYNTHESIZED_WIRE_712),
	.1GN(SYNTHESIZED_WIRE_713),
	.2A3(SYNTHESIZED_WIRE_500),
	.2GN(SYNTHESIZED_WIRE_713),
	.2A1(SYNTHESIZED_WIRE_712),
	.2A4(SYNTHESIZED_WIRE_503),
	.2A2(SYNTHESIZED_WIRE_712),
	.1Y2(Z80_LOCAL_DI[6]),
	.1Y4(Z80_LOCAL_DI[4]),
	.2Y1(Z80_LOCAL_DI[3]),
	.1Y1(Z80_LOCAL_DI[7]),
	.2Y3(Z80_LOCAL_DI[1]),
	.2Y4(Z80_LOCAL_DI[0]),
	.1Y3(Z80_LOCAL_DI[5]),
	.2Y2(Z80_LOCAL_DI[2]));

assign	SYNTHESIZED_WIRE_709 = OUT_pDBIN & SYNTHESIZED_WIRE_505;

assign	SYNTHESIZED_WIRE_710 = OUT_pDBIN & SYNTHESIZED_WIRE_506;

assign	SYNTHESIZED_WIRE_713 =  ~SYNTHESIZED_WIRE_710;


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_710 or SYNTHESIZED_WIRE_714)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_500 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SYNTHESIZED_WIRE_500 <= 1'b1;
else if (SYNTHESIZED_WIRE_710)
	SYNTHESIZED_WIRE_500 <= SYNTHESIZED_WIRE_714;
end



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_511 or Z80_LOCAL_D0[0])
begin
if (~IN_BOARD_RESET-)
		SPI_SD_CLK_SPEED <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		SPI_SD_CLK_SPEED <= 1'b1;
else if (SYNTHESIZED_WIRE_511)
	SPI_SD_CLK_SPEED <= Z80_LOCAL_D0;
end


\21mux 	b2v_inst479(
	.S(SPI_SD_CLK_SPEED),
	.B(400_KHz_CLK),
	.A(10mHz),
	.Y(LOCAL_SD_SPI_CLK));


\74138 	b2v_inst48(
	.A(S100_A0),
	.B(S100_A1),
	.G1(SYNTHESIZED_WIRE_513),
	.C(S100_A2),
	.G2AN(SYNTHESIZED_WIRE_716),
	.G2BN(SYNTHESIZED_WIRE_716),
	.Y0N(PORT_C0H-),
	.Y1N(PORT_C1H-),
	.Y2N(PORT_C2H-),
	
	
	
	.Y6N(PORT_C6H-),
	.Y7N(PORT_C7H-));


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_710 or SYNTHESIZED_WIRE_717)
begin
if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_503 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SYNTHESIZED_WIRE_503 <= 1'b1;
else if (SYNTHESIZED_WIRE_710)
	SYNTHESIZED_WIRE_503 <= SYNTHESIZED_WIRE_717;
end



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[7])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_7 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_7 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_7 <= DATA_FROM_SDCARD;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[6])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_6 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_6 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_6 <= DATA_FROM_SDCARD;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[5])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_5 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_5 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_5 <= DATA_FROM_SDCARD;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[4])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_4 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_4 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_4 <= DATA_FROM_SDCARD;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[3])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_3 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_3 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_3 <= DATA_FROM_SDCARD;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[2])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_2 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_2 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_2 <= DATA_FROM_SDCARD;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[1])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_1 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_1 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_1 <= DATA_FROM_SDCARD;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_711 or SYNTHESIZED_WIRE_709 or DATA_FROM_SDCARD[0])
begin
if (~IN_BOARD_RESET-)
		SDCARD_OUT_0 <= 1'b0;
else if (~SYNTHESIZED_WIRE_711)
		SDCARD_OUT_0 <= 1'b1;
else if (SYNTHESIZED_WIRE_709)
	SDCARD_OUT_0 <= DATA_FROM_SDCARD;
end

assign	SYNTHESIZED_WIRE_605 =  ~IN_BOARD_RESET-;


spi_master	b2v_inst490(
	.clock(LOCAL_SD_SPI_CLK),
	.reset_n(IN_BOARD_RESET-),
	.enable(SYNTHESIZED_WIRE_535),
	.cpol(SYNTHESIZED_WIRE_718),
	.cpha(SYNTHESIZED_WIRE_718),
	.cont(SYNTHESIZED_WIRE_718),
	.miso(SD_DO),
	.addr(SD_CARD_ADDRESS),
	.clk_div(SD_CARD_CLK_DIV),
	.tx_data(DATA_TO_SDCARD),
	.sclk(SD_CLK),
	.mosi(SD_CMD),
	.busy(SD_CARD_BUSY),
	.rx_data(DATA_FROM_SDCARD),
	.ss_n(SD_SLAVES));
	defparam	b2v_inst490.d_width = 8;
	defparam	b2v_inst490.slaves = 2;

assign	SYNTHESIZED_WIRE_505 =  ~PORT_SELECT_6C-;

assign	SYNTHESIZED_WIRE_506 =  ~PORT_SELECT_6E-;

assign	SYNTHESIZED_WIRE_708 =  ~SYNTHESIZED_WIRE_709;



always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[7])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[6])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[5])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[4])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[3])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


Counter01_32	b2v_inst5(
	.clock(2mHz),
	.q(COUNTER_BUS));

assign	OUT_RAM_READ- = ~(MEM_READ & SYNTHESIZED_WIRE_720);


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[2])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[1])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


always@(IN_BOARD_RESET- or SYNTHESIZED_WIRE_715 or SYNTHESIZED_WIRE_719 or Z80_LOCAL_D0[0])
begin
if (~IN_BOARD_RESET-)
		DATA_TO_SDCARD <= 1'b0;
else if (~SYNTHESIZED_WIRE_715)
		DATA_TO_SDCARD <= 1'b1;
else if (SYNTHESIZED_WIRE_719)
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
end


assign	SYNTHESIZED_WIRE_535 = SD_READ | SD_WRITE;



always@(posedge LOCAL_SD_SPI_CLK or negedge SYNTHESIZED_WIRE_706 or negedge SYNTHESIZED_WIRE_707)
begin
if (!SYNTHESIZED_WIRE_706)
	begin
	SD_WRITE <= 0;
	end
else
if (!SYNTHESIZED_WIRE_707)
	begin
	SD_WRITE <= 1;
	end
else
	begin
	SD_WRITE <= DFF_inst468;
	end
end

assign	SYNTHESIZED_WIRE_706 = SYNTHESIZED_WIRE_559 & IN_BOARD_RESET-;


always@(SYNTHESIZED_WIRE_715 or IN_BOARD_RESET- or SYNTHESIZED_WIRE_721 or Z80_LOCAL_D0[0])
begin
if (~SYNTHESIZED_WIRE_715)
		SYNTHESIZED_WIRE_714 <= 1'b0;
else if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_714 <= 1'b1;
else if (SYNTHESIZED_WIRE_721)
	SYNTHESIZED_WIRE_714 <= Z80_LOCAL_D0;
end


always@(SYNTHESIZED_WIRE_715 or IN_BOARD_RESET- or SYNTHESIZED_WIRE_721 or Z80_LOCAL_D0[1])
begin
if (~SYNTHESIZED_WIRE_715)
		SYNTHESIZED_WIRE_717 <= 1'b0;
else if (~IN_BOARD_RESET-)
		SYNTHESIZED_WIRE_717 <= 1'b1;
else if (SYNTHESIZED_WIRE_721)
	SYNTHESIZED_WIRE_717 <= Z80_LOCAL_D0;
end

assign	Z80_LOCAL_DI[1] = READ_RAM ? FPGA_BI_D1 : 1'bz;

assign	LED_1 = SD_SLAVES[0] | SD_SLAVES[0];

assign	SYNTHESIZED_WIRE_575 =  ~OUT_pDBIN;


always@(posedge SYNTHESIZED_WIRE_565 or negedge SYNTHESIZED_WIRE_722 or negedge SYNTHESIZED_WIRE_723)
begin
if (!SYNTHESIZED_WIRE_722)
	begin
	DFF_inst512 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_723)
	begin
	DFF_inst512 <= 1;
	end
else
	begin
	DFF_inst512 <= SYNTHESIZED_WIRE_723;
	end
end

assign	ROM_ADDRESS[13] = ROM_A13 | ROM_A13;


always@(posedge SYNTHESIZED_WIRE_568 or negedge IN_BOARD_RESET- or negedge SYNTHESIZED_WIRE_569)
begin
if (!IN_BOARD_RESET-)
	begin
	ROM_A13 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_569)
	begin
	ROM_A13 <= 1;
	end
else
	begin
	ROM_A13 <= Z80_LOCAL_D0[2];
	end
end




always@(posedge LOCAL_SD_SPI_CLK or negedge SYNTHESIZED_WIRE_722 or negedge SYNTHESIZED_WIRE_723)
begin
if (!SYNTHESIZED_WIRE_722)
	begin
	SD_READ <= 0;
	end
else
if (!SYNTHESIZED_WIRE_723)
	begin
	SD_READ <= 1;
	end
else
	begin
	SD_READ <= DFF_inst512;
	end
end

assign	SD_CARD_CLK_DIV =  ~SYNTHESIZED_WIRE_724;


assign	USB_DATA_IN- =  ~USB_DATA_IN;

assign	SD_CARD_ADDRESS =  ~SYNTHESIZED_WIRE_724;

assign	SYNTHESIZED_WIRE_574 =  ~SD_CARD_BUSY;

assign	SYNTHESIZED_WIRE_722 = SYNTHESIZED_WIRE_574 & IN_BOARD_RESET-;

assign	SYNTHESIZED_WIRE_486 = ~(PORT_SELECT_6F- | OUT_pWR-);

assign	SYNTHESIZED_WIRE_565 = ~(PORT_SELECT_6F- | SYNTHESIZED_WIRE_575);

assign	SYNTHESIZED_WIRE_559 =  ~SD_CARD_BUSY;

assign	SYNTHESIZED_WIRE_576 =  ~OUT_sOUT;

assign	SYNTHESIZED_WIRE_90 = SD_CARD_READ_DATA- & USB_STATUS_IN- & USB_DATA_IN-;

assign	SYNTHESIZED_WIRE_568 = ~(SYNTHESIZED_WIRE_576 | OUT_pWR- | PORT_7-);

assign	SYNTHESIZED_WIRE_675 = ROM_A13 | ROM_A12;


\74157 	b2v_inst53(
	.A1(SYNTHESIZED_WIRE_577),
	.B1(SYNTHESIZED_WIRE_725),
	.SEL(SYNTHESIZED_WIRE_638),
	.B2(SYNTHESIZED_WIRE_725),
	.A3(SYNTHESIZED_WIRE_581),
	.B3(SYNTHESIZED_WIRE_725),
	.A2(SYNTHESIZED_WIRE_583),
	.B4(SYNTHESIZED_WIRE_725),
	.GN(SYNTHESIZED_WIRE_725),
	.A4(SYNTHESIZED_WIRE_586),
	.Y2(S100_A9),
	.Y1(S100_A8),
	.Y4(S100_A11),
	.Y3(S100_A10));

assign	SYNTHESIZED_WIRE_91 = BAR_IN_ENABLE- & SYNTHESIZED_WIRE_587 & SYNTHESIZED_WIRE_588;

assign	SYNTHESIZED_WIRE_587 =  ~PS2_STATUS_IN;

assign	SYNTHESIZED_WIRE_588 =  ~PS2_DATA_IN;


assign	IO_OUTPUT = Z80_WR & Z80_IORQ;

assign	IO_INPUT = Z80_IORQ & Z80_RD;

assign	MEM_READ = Z80_RD & Z80_MREQ;

assign	SYNTHESIZED_WIRE_726 = Z80_MREQ & Z80_RFSH-;


\74373 	b2v_inst59(
	.D1(SYNTHESIZED_WIRE_589),
	.D3(IO_INPUT),
	.D6(Z80_M1),
	.D7(Z80_INTA),
	.D2(IO_OUTPUT),
	.G(ADDRESS_LATCH),
	.D4(MEM_READ),
	.D5(SYNTHESIZED_WIRE_590),
	
	.OEN(SYNTHESIZED_WIRE_591),
	.Q3(OUT_sINP),
	.Q6(OUT_sM1),
	.Q7(OUT_sINTA),
	.Q2(OUT_sOUT),
	
	.Q4(OUT_sMEMR),
	.Q5(OUT_sWO-),
	.Q1(OUT_sHLTA));

assign	IOBYTE_OE- = IOBYTE- | SYNTHESIZED_WIRE_640;

assign	SYNTHESIZED_WIRE_595 = ~(Z80_RD- & SYNTHESIZED_WIRE_726);

assign	SYNTHESIZED_WIRE_670 = ~(Z80_IORQ & Z80_M1);

assign	SYNTHESIZED_WIRE_665 =  ~OUT_pDBIN;

assign	MEM_WRITE = Z80_WR & Z80_MREQ;


assign	Z80_INTA =  ~SYNTHESIZED_WIRE_670;

assign	OUT_CPU_CLK- =  ~OUT_CPU_CLK;


assign	WRITE = ~(Z80_WR- & SYNTHESIZED_WIRE_595);

assign	SYNTHESIZED_WIRE_590 =  ~WRITE;


vga80x40	b2v_inst7(
	.reset(IN_BOARD_RESET),
	.clk25MHz(25Mhz),
	.FONT_D(FONT_D),
	.ocrx(ocrx),
	.ocry(ocry),
	.octl(CTL),
	.TEXT_D(RAM_TEXT_D),
	.R(VGA_R),
	.G(VGA_G),
	.B(VGA_B),
	.hsync(HSync),
	.vsync(VSync),
	.cursor_x(CURSOR_X[6:0]),
	.cursor_y(CURSOR_Y[5:0]),
	.FONT_A(FONT_A),
	.TEXT_A(TEXT_A));

assign	START_SYNC = ~(Z80_INTA | SYNTHESIZED_WIRE_726 | DFF_inst92);


\74244 	b2v_inst71(
	.1A2(pSYNC_RAW),
	.1A4(SYNTHESIZED_WIRE_727),
	.1A1(DFF_inst97),
	.1A3(ADDRESS_LATCH),
	.1GN(SYNTHESIZED_WIRE_598),
	.2A3(SYNTHESIZED_WIRE_599),
	.2GN(SYNTHESIZED_WIRE_600),
	.2A1(OUT_CPU_CLK),
	.2A4(FPGA_IN_INT-),
	.2A2(2mHz),
	.1Y2(FPGA_OUT_pSYNC),
	.1Y4(OUT_pWR-),
	.2Y1(FPGA_OUT_PHI),
	.1Y1(OUT_pDBIN),
	.2Y3(OUT_MWRT),
	.2Y4(S100_INT-),
	.1Y3(FPGA_OUT_pSTVAL-),
	.2Y2(FPGA_OUT_2mHz_CLOCK));

assign	SYNTHESIZED_WIRE_613 =  ~START_SYNC;

assign	JMP_ENABLE =  ~JMP_ENABLE-;

assign	OUT_RAM_WRITE- = ~(MEM_WRITE & SYNTHESIZED_WIRE_720);



assign	SYNTHESIZED_WIRE_666 = PORT_C0H- | SYNTHESIZED_WIRE_665;

assign	SYNTHESIZED_WIRE_32 =  ~SYNTHESIZED_WIRE_603;

assign	Z80_LOCAL_DI[7] = ROM_OE ? SYNTHESIZED_WIRE_604[7] : 1'bz;
assign	Z80_LOCAL_DI[6] = ROM_OE ? SYNTHESIZED_WIRE_604[6] : 1'bz;
assign	Z80_LOCAL_DI[5] = ROM_OE ? SYNTHESIZED_WIRE_604[5] : 1'bz;
assign	Z80_LOCAL_DI[4] = ROM_OE ? SYNTHESIZED_WIRE_604[4] : 1'bz;
assign	Z80_LOCAL_DI[3] = ROM_OE ? SYNTHESIZED_WIRE_604[3] : 1'bz;
assign	Z80_LOCAL_DI[2] = ROM_OE ? SYNTHESIZED_WIRE_604[2] : 1'bz;
assign	Z80_LOCAL_DI[1] = ROM_OE ? SYNTHESIZED_WIRE_604[1] : 1'bz;
assign	Z80_LOCAL_DI[0] = ROM_OE ? SYNTHESIZED_WIRE_604[0] : 1'bz;


uart	b2v_inst8(
	.clk(50mHz),
	.rst(SYNTHESIZED_WIRE_605),
	.rx(DATA_FROM_USB_PORT),
	.transmit(SYNTHESIZED_WIRE_606),
	.data_read(USB_DATA_IN),
	.tx_byte(USB_DATA_OUT_BUS),
	.tx(SERIAL_DATA_TO_USB_PORT),
	.received(UART_Byte_Recieved),
	.is_receiving(UART_Busy_Recieving),
	.is_transmitting(UART_Busy_Transmitting),
	.recv_error(UART_Error),
	.data_ready(UART_DATA_READY),
	.rx_byte(USB_DATA_IN_BUS));
	defparam	b2v_inst8.CLOCK_DIVIDE = 1303;
	defparam	b2v_inst8.FLAG_HIGH = 1;
	defparam	b2v_inst8.FLAG_LOW = 0;
	defparam	b2v_inst8.RX_CHECK_START = 1;
	defparam	b2v_inst8.RX_CHECK_STOP = 3;
	defparam	b2v_inst8.RX_DELAY_RESTART = 4;
	defparam	b2v_inst8.RX_ERROR = 5;
	defparam	b2v_inst8.RX_IDLE = 0;
	defparam	b2v_inst8.RX_READ_BITS = 2;
	defparam	b2v_inst8.RX_RECEIVED = 6;
	defparam	b2v_inst8.TX_DELAY_RESTART = 2;
	defparam	b2v_inst8.TX_IDLE = 0;
	defparam	b2v_inst8.TX_SENDING = 1;

assign	END_SYNC =  ~DFF_inst95;

assign	SYNTHESIZED_WIRE_727 = ~(Z80_WR & END_SYNC);


assign	SYNTHESIZED_WIRE_599 = ~(SYNTHESIZED_WIRE_727 | IO_OUTPUT);

assign	SYNTHESIZED_WIRE_600 =  ~SYNTHESIZED_WIRE_681;

assign	SYNTHESIZED_WIRE_603 =  ~ADDRESS_LATCH;

assign	SYNTHESIZED_WIRE_598 =  ~IN_CDSB-;

assign	FPGA_OUT_CTL_OE- =  ~IN_CDSB-;

assign	FPGA_OUT_STATUS_OE- =  ~IN_SDSB-;


assign	FPGA_OUT_LOW_ROM_LED- = SYNTHESIZED_WIRE_675 | DISABLE_ALL_ROM;




always@(posedge OUT_CPU_CLK or negedge Z80_IORQ or negedge SYNTHESIZED_WIRE_609)
begin
if (!Z80_IORQ)
	begin
	DFF_inst92 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_609)
	begin
	DFF_inst92 <= 1;
	end
else
	begin
	DFF_inst92 <= Z80_IORQ;
	end
end


always@(posedge OUT_CPU_CLK or negedge SYNTHESIZED_WIRE_728 or negedge IN_BOARD_RESET-)
begin
if (!SYNTHESIZED_WIRE_728)
	begin
	SYNTHESIZED_WIRE_681 <= 0;
	end
else
if (!IN_BOARD_RESET-)
	begin
	SYNTHESIZED_WIRE_681 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_681 <= SYNTHESIZED_WIRE_728;
	end
end



always@(posedge OUT_CPU_CLK or negedge SYNTHESIZED_WIRE_612 or negedge SYNTHESIZED_WIRE_613)
begin
if (!SYNTHESIZED_WIRE_612)
	begin
	DFF_inst95 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_613)
	begin
	DFF_inst95 <= 1;
	end
else
	begin
	DFF_inst95 <= START_SYNC;
	end
end



always@(posedge SYNTHESIZED_WIRE_615 or negedge SYNTHESIZED_WIRE_729 or negedge SYNTHESIZED_WIRE_617)
begin
if (!SYNTHESIZED_WIRE_729)
	begin
	DFF_inst97 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_617)
	begin
	DFF_inst97 <= 1;
	end
else
	begin
	DFF_inst97 <= SYNTHESIZED_WIRE_729;
	end
end


assign	FPGA_OUT_RAM_OE- = OUT_RAM_READ- & OUT_RAM_WRITE-;

assign	FPGA_OUT_A1 = S100_A1;
assign	IN_BOARD_RESET- = FPGA_IN_BOARD_RESET-;
assign	DIP_7 = DIP0;
assign	IN_SDSB- = FPGA_IN_SDSB-;
assign	IN_CDSB- = FPGA_IN_CDSB-;
assign	50mHz = CLK_50;
assign	DATA_FROM_USB_PORT = USB_RX;
assign	DIP_5 = DIP2;
assign	DIP_6 = DIP1;
assign	FPGA_OUT_A2 = S100_A2;
assign	FPGA_OUT_A3 = S100_A3;
assign	FPGA_OUT_A4 = S100_A4;
assign	FPGA_OUT_A5 = S100_A5;
assign	FPGA_OUT_A6 = S100_A6;
assign	FPGA_OUT_A7 = S100_A7;
assign	FPGA_OUT_A16 = S100_A16;
assign	FPGA_OUT_A17 = S100_A17;
assign	FPGA_OUT_A18 = S100_A18;
assign	FPGA_OUT_A19 = S100_A19;
assign	FPGA_OUT_CPU_CLK = OUT_CPU_CLK-;
assign	FPGA_OUT_sINTA = OUT_sINTA;
assign	FPGA_OUT_sM1 = OUT_sM1;
assign	FPGA_OUT_sWO- = OUT_sWO-;
assign	FPGA_OUT_sMEMR = OUT_sMEMR;
assign	FPGA_OUT_sINP = OUT_sINP;
assign	FPGA_OUT_sOUT = OUT_sOUT;
assign	FPGA_OUT_sHLTA = OUT_sHLTA;
assign	FPGA_OUT_pDBIN = OUT_pDBIN;
assign	FPGA_OUT_pWR- = OUT_pWR-;
assign	FPGA_OUT_MWRT = OUT_MWRT;
assign	FPGA_OUT_RAM_WR- = OUT_RAM_WRITE-;
assign	FPGA_OUT_DO0 = DATA_OUT_D0;
assign	FPGA_OUT_DO1 = DATA_OUT_D1;
assign	FPGA_OUT_DO2 = DATA_OUT_D2;
assign	FPGA_OUT_DO3 = DATA_OUT_D3;
assign	FPGA_OUT_DO4 = DATA_OUT_D4;
assign	FPGA_OUT_DO5 = DATA_OUT_D5;
assign	FPGA_OUT_DO6 = DATA_OUT_D6;
assign	FPGA_OUT_DO7 = DATA_OUT_D7;
assign	FPGA_OUT_A0 = S100_A0;
assign	FPGA_OUT_A8 = S100_A8;
assign	FPGA_OUT_A9 = S100_A9;
assign	FPGA_OUT_A11 = S100_A11;
assign	FPGA_OUT_A10 = S100_A10;
assign	FPGA_OUT_A12 = S100_A12;
assign	FPGA_OUT_A13 = S100_A13;
assign	FPGA_OUT_A14 = S100_A14;
assign	FPGA_OUT_A15 = S100_A15;
assign	USB_TX = SERIAL_DATA_TO_USB_PORT;
assign	RTC_SPI_CLK = SPI_MASTER_CLK;
assign	DIAG_LED = SPI_SD_CLK_SPEED;
assign	FPGA_OUT_SPARE1 = LOCAL_SD_SPI_CLK;

endmodule
