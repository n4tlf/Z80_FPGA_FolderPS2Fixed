-- Copyright (C) 2021  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 21.1.0 Build 842 10/21/2021 SJ Lite Edition"
-- CREATED		"Thu Mar 31 16:17:06 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Z80_FPGA IS 
	PORT
	(
		CLK_50 :  IN  STD_LOGIC;
		FPGA_IN_XRDY :  IN  STD_LOGIC;
		FPGA_IN_RDY :  IN  STD_LOGIC;
		FPGA_IN_SDSB- :  IN  STD_LOGIC;
		FPGA_IN_CDSB- :  IN  STD_LOGIC;
		FPGA_IN_pHOLD- :  IN  STD_LOGIC;
		FPGA_IN_DI0 :  IN  STD_LOGIC;
		FPGA_IN_DI1 :  IN  STD_LOGIC;
		FPGA_IN_DI2 :  IN  STD_LOGIC;
		FPGA_IN_DI4 :  IN  STD_LOGIC;
		FPGA_IN_DI5 :  IN  STD_LOGIC;
		FPGA_IN_DI6 :  IN  STD_LOGIC;
		FPGA_IN_DI7 :  IN  STD_LOGIC;
		FPGA_IN_DI3 :  IN  STD_LOGIC;
		FPGA_IN_PS2_CLK :  IN  STD_LOGIC;
		FPGA_IN_PS2_DATA :  IN  STD_LOGIC;
		FPGA_IN_PRN_ACK :  IN  STD_LOGIC;
		FPGA_IN_PRN_BUSY :  IN  STD_LOGIC;
		RTC_SPI_SO :  IN  STD_LOGIC;
		DIP7 :  IN  STD_LOGIC;
		DIP6 :  IN  STD_LOGIC;
		DIP5 :  IN  STD_LOGIC;
		DIP4 :  IN  STD_LOGIC;
		DIP3 :  IN  STD_LOGIC;
		DIP2 :  IN  STD_LOGIC;
		DIP1 :  IN  STD_LOGIC;
		DIP0 :  IN  STD_LOGIC;
		FPGA_IN_INT_B- :  IN  STD_LOGIC;
		FPGA_IN_INT_C- :  IN  STD_LOGIC;
		FPGA_IN_INT_D- :  IN  STD_LOGIC;
		FPGA_IN_INT_A- :  IN  STD_LOGIC;
		USB_RX :  IN  STD_LOGIC;
		FPGA_IN_INT- :  IN  STD_LOGIC;
		RTC_INT :  IN  STD_LOGIC;
		FPGA_IN_ENABLE_INTA :  IN  STD_LOGIC;
		FPGA_IN_BOARD_RESET- :  IN  STD_LOGIC;
		SD_DO :  IN  STD_LOGIC;
		FPGA_BI_D0 :  INOUT  STD_LOGIC;
		FPGA_BI_D1 :  INOUT  STD_LOGIC;
		FPGA_BI_D2 :  INOUT  STD_LOGIC;
		FPGA_BI_D3 :  INOUT  STD_LOGIC;
		FPGA_BI_D4 :  INOUT  STD_LOGIC;
		FPGA_BI_D5 :  INOUT  STD_LOGIC;
		FPGA_BI_D6 :  INOUT  STD_LOGIC;
		FPGA_BI_D7 :  INOUT  STD_LOGIC;
		FPGA_OUT_A1 :  OUT  STD_LOGIC;
		FPGA_OUT_A2 :  OUT  STD_LOGIC;
		FPGA_OUT_A3 :  OUT  STD_LOGIC;
		FPGA_OUT_A4 :  OUT  STD_LOGIC;
		FPGA_OUT_A5 :  OUT  STD_LOGIC;
		FPGA_OUT_A6 :  OUT  STD_LOGIC;
		FPGA_OUT_A7 :  OUT  STD_LOGIC;
		FPGA_OUT_A16 :  OUT  STD_LOGIC;
		FPGA_OUT_A17 :  OUT  STD_LOGIC;
		FPGA_OUT_A18 :  OUT  STD_LOGIC;
		FPGA_OUT_A19 :  OUT  STD_LOGIC;
		FPGA_OUT_CPU_CLK :  OUT  STD_LOGIC;
		FPGA_OUT_sINTA :  OUT  STD_LOGIC;
		FPGA_OUT_sM1 :  OUT  STD_LOGIC;
		FPGA_OUT_sWO- :  OUT  STD_LOGIC;
		FPGA_OUT_sMEMR :  OUT  STD_LOGIC;
		FPGA_OUT_sINP :  OUT  STD_LOGIC;
		FPGA_OUT_sOUT :  OUT  STD_LOGIC;
		FPGA_OUT_sHLTA :  OUT  STD_LOGIC;
		FPGA_OUT_pDBIN :  OUT  STD_LOGIC;
		FPGA_OUT_pWR- :  OUT  STD_LOGIC;
		FPGA_OUT_MWRT :  OUT  STD_LOGIC;
		FPGA_OUT_2mHz_CLOCK :  OUT  STD_LOGIC;
		FPGA_OUT_PHI :  OUT  STD_LOGIC;
		FPGA_OUT_pSYNC :  OUT  STD_LOGIC;
		FPGA_OUT_pSTVAL- :  OUT  STD_LOGIC;
		FPGA_OUT_RAM_WR- :  OUT  STD_LOGIC;
		FPGA_OUT_RAM_OE- :  OUT  STD_LOGIC;
		FPGA_OUT_DO0 :  OUT  STD_LOGIC;
		FPGA_OUT_DO1 :  OUT  STD_LOGIC;
		FPGA_OUT_DO2 :  OUT  STD_LOGIC;
		FPGA_OUT_DO3 :  OUT  STD_LOGIC;
		FPGA_OUT_DO4 :  OUT  STD_LOGIC;
		FPGA_OUT_DO5 :  OUT  STD_LOGIC;
		FPGA_OUT_DO6 :  OUT  STD_LOGIC;
		FPGA_OUT_DO7 :  OUT  STD_LOGIC;
		FPGA_OUT_A0 :  OUT  STD_LOGIC;
		FPGA_OUT_A8 :  OUT  STD_LOGIC;
		FPGA_OUT_A9 :  OUT  STD_LOGIC;
		FPGA_OUT_A11 :  OUT  STD_LOGIC;
		FPGA_OUT_A10 :  OUT  STD_LOGIC;
		FPGA_OUT_A12 :  OUT  STD_LOGIC;
		FPGA_OUT_A13 :  OUT  STD_LOGIC;
		FPGA_OUT_A14 :  OUT  STD_LOGIC;
		FPGA_OUT_A15 :  OUT  STD_LOGIC;
		FPGA_OUT_STATUS_DISABLE :  OUT  STD_LOGIC;
		FPGA_OUT_pHLDA :  OUT  STD_LOGIC;
		FPGA_OUT_CTL_DISABLE :  OUT  STD_LOGIC;
		FPGA_OUT_CTL_OE- :  OUT  STD_LOGIC;
		FPGA_OUT_STATUS_OE- :  OUT  STD_LOGIC;
		FPGA_ADD_OE- :  OUT  STD_LOGIC;
		FPGA_OUT_DO_OE- :  OUT  STD_LOGIC;
		FPGA_OUT_DI_OE- :  OUT  STD_LOGIC;
		FPGA_OUT_RAM_CS- :  OUT  STD_LOGIC;
		FPGA_OUT_RAM_A17 :  OUT  STD_LOGIC;
		FPGA_OUT_RAM_A18 :  OUT  STD_LOGIC;
		FPGA_OUT_RAM_A16 :  OUT  STD_LOGIC;
		USB_TX :  OUT  STD_LOGIC;
		F_BAR0 :  OUT  STD_LOGIC;
		F_BAR1 :  OUT  STD_LOGIC;
		F_BAR2 :  OUT  STD_LOGIC;
		F_BAR3 :  OUT  STD_LOGIC;
		F_BAR4 :  OUT  STD_LOGIC;
		F_BAR5 :  OUT  STD_LOGIC;
		F_BAR6 :  OUT  STD_LOGIC;
		F_BAR7 :  OUT  STD_LOGIC;
		USB_TX_BUSY_LED :  OUT  STD_LOGIC;
		USB_RX_BUSY_LED :  OUT  STD_LOGIC;
		5V_OUT_IDE_PORTS_RD- :  OUT  STD_LOGIC;
		5V_OUT_IDE_PORTS_WR- :  OUT  STD_LOGIC;
		VGA_R :  OUT  STD_LOGIC;
		VGA_G :  OUT  STD_LOGIC;
		VGA_B :  OUT  STD_LOGIC;
		HSync :  OUT  STD_LOGIC;
		VSync :  OUT  STD_LOGIC;
		BUZZER :  OUT  STD_LOGIC;
		F_BOARD_ACTIVE- :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_0 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_1 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_2 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_3 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_4 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_5 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_6 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_7 :  OUT  STD_LOGIC;
		FPGA_OUT_PRN_STROBE :  OUT  STD_LOGIC;
		PRN_ACK_LED :  OUT  STD_LOGIC;
		FPGA_OUT_PHANTOM :  OUT  STD_LOGIC;
		S100_PHANTOM_LED :  OUT  STD_LOGIC;
		RTC_CS :  OUT  STD_LOGIC;
		RTC_SPI_SI :  OUT  STD_LOGIC;
		RTC_SPI_CLK :  OUT  STD_LOGIC;
		SD_CMD :  OUT  STD_LOGIC;
		SD_CLK :  OUT  STD_LOGIC;
		LED_4 :  OUT  STD_LOGIC;
		P1 :  OUT  STD_LOGIC;
		LED_1 :  OUT  STD_LOGIC;
		DIAG_LED :  OUT  STD_LOGIC;
		SD_CS_B- :  OUT  STD_LOGIC;
		FPGA_OUT_SPARE1 :  OUT  STD_LOGIC;
		SD_CS_A- :  OUT  STD_LOGIC;
		FPGA_OUT_IDE_RD- :  OUT  STD_LOGIC;
		FPGA_OUT_IDE_WR- :  OUT  STD_LOGIC;
		FPGA_OUT_8255_SEL- :  OUT  STD_LOGIC;
		FPGA_OUT_HIGH_ROM_LED- :  OUT  STD_LOGIC;
		FPGA_OUT_LOW_ROM_LED- :  OUT  STD_LOGIC;
		FPGA_OUT_HIGH_RAM_LED- :  OUT  STD_LOGIC;
		LED_2 :  OUT  STD_LOGIC;
		LED_3 :  OUT  STD_LOGIC
	);
END Z80_FPGA;

ARCHITECTURE bdf_type OF Z80_FPGA IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT \21mux_19\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_19\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_19\: COMPONENT IS true;

COMPONENT \21mux_35\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_35\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_35\: COMPONENT IS true;

COMPONENT \74138_11\
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 G1 : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 G2AN : IN STD_LOGIC;
		 G2BN : IN STD_LOGIC;
		 Y0N : OUT STD_LOGIC;
		 Y2N : OUT STD_LOGIC;
		 Y3N : OUT STD_LOGIC;
		 Y6N : OUT STD_LOGIC;
		 Y7N : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74138_11\: COMPONENT IS true;
ATTRIBUTE noopt OF \74138_11\: COMPONENT IS true;

COMPONENT \74138_22\
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 G1 : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 G2AN : IN STD_LOGIC;
		 G2BN : IN STD_LOGIC;
		 Y0N : OUT STD_LOGIC;
		 Y1N : OUT STD_LOGIC;
		 Y2N : OUT STD_LOGIC;
		 Y3N : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74138_22\: COMPONENT IS true;
ATTRIBUTE noopt OF \74138_22\: COMPONENT IS true;

COMPONENT \74138_27\
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 G1 : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 G2AN : IN STD_LOGIC;
		 G2BN : IN STD_LOGIC;
		 Y0N : OUT STD_LOGIC;
		 Y1N : OUT STD_LOGIC;
		 Y2N : OUT STD_LOGIC;
		 Y3N : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74138_27\: COMPONENT IS true;
ATTRIBUTE noopt OF \74138_27\: COMPONENT IS true;

COMPONENT \74138_36\
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 G1 : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 G2AN : IN STD_LOGIC;
		 G2BN : IN STD_LOGIC;
		 Y0N : OUT STD_LOGIC;
		 Y1N : OUT STD_LOGIC;
		 Y2N : OUT STD_LOGIC;
		 Y6N : OUT STD_LOGIC;
		 Y7N : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74138_36\: COMPONENT IS true;
ATTRIBUTE noopt OF \74138_36\: COMPONENT IS true;

COMPONENT \74138_7\
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 G1 : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 G2AN : IN STD_LOGIC;
		 G2BN : IN STD_LOGIC;
		 Y0N : OUT STD_LOGIC;
		 Y1N : OUT STD_LOGIC;
		 Y2N : OUT STD_LOGIC;
		 Y3N : OUT STD_LOGIC;
		 Y4N : OUT STD_LOGIC;
		 Y5N : OUT STD_LOGIC;
		 Y6N : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74138_7\: COMPONENT IS true;
ATTRIBUTE noopt OF \74138_7\: COMPONENT IS true;

COMPONENT \74148_25\
	PORT(5N : IN STD_LOGIC;
		 0N : IN STD_LOGIC;
		 1N : IN STD_LOGIC;
		 2N : IN STD_LOGIC;
		 3N : IN STD_LOGIC;
		 4N : IN STD_LOGIC;
		 EIN : IN STD_LOGIC;
		 6N : IN STD_LOGIC;
		 7N : IN STD_LOGIC;
		 A1N : OUT STD_LOGIC;
		 A0N : OUT STD_LOGIC;
		 A2N : OUT STD_LOGIC;
		 GSN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74148_25\: COMPONENT IS true;
ATTRIBUTE noopt OF \74148_25\: COMPONENT IS true;

COMPONENT \74157_37\
	PORT(A1 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 SEL : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 GN : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 Y2 : OUT STD_LOGIC;
		 Y1 : OUT STD_LOGIC;
		 Y4 : OUT STD_LOGIC;
		 Y3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74157_37\: COMPONENT IS true;
ATTRIBUTE noopt OF \74157_37\: COMPONENT IS true;

COMPONENT \74157_8\
	PORT(A1 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 SEL : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 A3 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 GN : IN STD_LOGIC;
		 A4 : IN STD_LOGIC;
		 Y2 : OUT STD_LOGIC;
		 Y1 : OUT STD_LOGIC;
		 Y4 : OUT STD_LOGIC;
		 Y3 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74157_8\: COMPONENT IS true;
ATTRIBUTE noopt OF \74157_8\: COMPONENT IS true;

COMPONENT \74164_24\
	PORT(CLRN : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 QB : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74164_24\: COMPONENT IS true;
ATTRIBUTE noopt OF \74164_24\: COMPONENT IS true;

COMPONENT \74165_0\
	PORT(D : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 H : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 CLKIH : IN STD_LOGIC;
		 E : IN STD_LOGIC;
		 F : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 STLD : IN STD_LOGIC;
		 SER : IN STD_LOGIC;
		 QHN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74165_0\: COMPONENT IS true;
ATTRIBUTE noopt OF \74165_0\: COMPONENT IS true;

COMPONENT \74165_4\
	PORT(D : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 H : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 CLKIH : IN STD_LOGIC;
		 E : IN STD_LOGIC;
		 F : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 STLD : IN STD_LOGIC;
		 SER : IN STD_LOGIC;
		 QHN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74165_4\: COMPONENT IS true;
ATTRIBUTE noopt OF \74165_4\: COMPONENT IS true;

COMPONENT \74244_13\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_13\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_13\: COMPONENT IS true;

COMPONENT \74244_14\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_14\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_14\: COMPONENT IS true;

COMPONENT \74244_23\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_23\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_23\: COMPONENT IS true;

COMPONENT \74244_29\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_29\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_29\: COMPONENT IS true;

COMPONENT \74244_31\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_31\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_31\: COMPONENT IS true;

COMPONENT \74244_32\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_32\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_32\: COMPONENT IS true;

COMPONENT \74244_33\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_33\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_33\: COMPONENT IS true;

COMPONENT \74244_34\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_34\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_34\: COMPONENT IS true;

COMPONENT \74244_39\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_39\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_39\: COMPONENT IS true;

COMPONENT \74373_1\
	PORT(D1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D6 : IN STD_LOGIC;
		 D7 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 D4 : IN STD_LOGIC;
		 D5 : IN STD_LOGIC;
		 D8 : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q6 : OUT STD_LOGIC;
		 Q7 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC;
		 Q8 : OUT STD_LOGIC;
		 Q4 : OUT STD_LOGIC;
		 Q5 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74373_1\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373_1\: COMPONENT IS true;

COMPONENT \74373_10\
	PORT(D1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D6 : IN STD_LOGIC;
		 D7 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 D4 : IN STD_LOGIC;
		 D5 : IN STD_LOGIC;
		 D8 : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q6 : OUT STD_LOGIC;
		 Q7 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC;
		 Q8 : OUT STD_LOGIC;
		 Q4 : OUT STD_LOGIC;
		 Q5 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74373_10\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373_10\: COMPONENT IS true;

COMPONENT \74373_2\
	PORT(D1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D6 : IN STD_LOGIC;
		 D7 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 D4 : IN STD_LOGIC;
		 D5 : IN STD_LOGIC;
		 D8 : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q6 : OUT STD_LOGIC;
		 Q7 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC;
		 Q8 : OUT STD_LOGIC;
		 Q4 : OUT STD_LOGIC;
		 Q5 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74373_2\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373_2\: COMPONENT IS true;

COMPONENT \74373_26\
	PORT(D1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D6 : IN STD_LOGIC;
		 D7 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 D4 : IN STD_LOGIC;
		 D5 : IN STD_LOGIC;
		 D8 : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q6 : OUT STD_LOGIC;
		 Q7 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC;
		 Q8 : OUT STD_LOGIC;
		 Q4 : OUT STD_LOGIC;
		 Q5 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74373_26\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373_26\: COMPONENT IS true;

COMPONENT \74373_3\
	PORT(D1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D6 : IN STD_LOGIC;
		 D7 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 D4 : IN STD_LOGIC;
		 D5 : IN STD_LOGIC;
		 D8 : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC;
		 Q4 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74373_3\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373_3\: COMPONENT IS true;

COMPONENT \74373_38\
	PORT(D1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D6 : IN STD_LOGIC;
		 D7 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 D4 : IN STD_LOGIC;
		 D5 : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 Q3 : OUT STD_LOGIC;
		 Q6 : OUT STD_LOGIC;
		 Q7 : OUT STD_LOGIC;
		 Q2 : OUT STD_LOGIC;
		 Q4 : OUT STD_LOGIC;
		 Q5 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74373_38\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373_38\: COMPONENT IS true;

COMPONENT \74373b_15\
	PORT(G : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(8 DOWNTO 1);
		 Q : OUT STD_LOGIC_VECTOR(8 DOWNTO 1));
END COMPONENT;
ATTRIBUTE black_box OF \74373b_15\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373b_15\: COMPONENT IS true;

COMPONENT \74373b_16\
	PORT(G : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(8 DOWNTO 1);
		 Q : OUT STD_LOGIC_VECTOR(8 DOWNTO 1));
END COMPONENT;
ATTRIBUTE black_box OF \74373b_16\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373b_16\: COMPONENT IS true;

COMPONENT \74373b_17\
	PORT(G : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(8 DOWNTO 1);
		 Q : OUT STD_LOGIC_VECTOR(8 DOWNTO 1));
END COMPONENT;
ATTRIBUTE black_box OF \74373b_17\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373b_17\: COMPONENT IS true;

COMPONENT \74373b_18\
	PORT(G : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(8 DOWNTO 1);
		 Q : OUT STD_LOGIC_VECTOR(8 DOWNTO 1));
END COMPONENT;
ATTRIBUTE black_box OF \74373b_18\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373b_18\: COMPONENT IS true;

COMPONENT \74373b_21\
	PORT(G : IN STD_LOGIC;
		 OEN : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(8 DOWNTO 1);
		 Q : OUT STD_LOGIC_VECTOR(8 DOWNTO 1));
END COMPONENT;
ATTRIBUTE black_box OF \74373b_21\: COMPONENT IS true;
ATTRIBUTE noopt OF \74373b_21\: COMPONENT IS true;

COMPONENT \74684_12\
	PORT(P2 : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 P1 : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 P0 : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 P7 : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 P6 : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 P5 : IN STD_LOGIC;
		 P4 : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 P3 : IN STD_LOGIC;
		 EQUALN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74684_12\: COMPONENT IS true;
ATTRIBUTE noopt OF \74684_12\: COMPONENT IS true;

COMPONENT \74684_20\
	PORT(P2 : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 P1 : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 P0 : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 P7 : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 P6 : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 P5 : IN STD_LOGIC;
		 P4 : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 P3 : IN STD_LOGIC;
		 EQUALN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74684_20\: COMPONENT IS true;
ATTRIBUTE noopt OF \74684_20\: COMPONENT IS true;

COMPONENT \74684_28\
	PORT(P2 : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 P1 : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 P0 : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 P7 : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 P6 : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 P5 : IN STD_LOGIC;
		 P4 : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 P3 : IN STD_LOGIC;
		 EQUALN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74684_28\: COMPONENT IS true;
ATTRIBUTE noopt OF \74684_28\: COMPONENT IS true;

COMPONENT \74684_30\
	PORT(P2 : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 P1 : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 P0 : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 P7 : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 P6 : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 P5 : IN STD_LOGIC;
		 P4 : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 P3 : IN STD_LOGIC;
		 EQUALN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74684_30\: COMPONENT IS true;
ATTRIBUTE noopt OF \74684_30\: COMPONENT IS true;

COMPONENT \74684_5\
	PORT(P2 : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 P1 : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 P0 : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 P7 : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 P6 : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 P5 : IN STD_LOGIC;
		 P4 : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 P3 : IN STD_LOGIC;
		 EQUALN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74684_5\: COMPONENT IS true;
ATTRIBUTE noopt OF \74684_5\: COMPONENT IS true;

COMPONENT \74684_6\
	PORT(P2 : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 P1 : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 P0 : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 P7 : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 P6 : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 P5 : IN STD_LOGIC;
		 P4 : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 P3 : IN STD_LOGIC;
		 EQUALN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74684_6\: COMPONENT IS true;
ATTRIBUTE noopt OF \74684_6\: COMPONENT IS true;

COMPONENT \74684_9\
	PORT(P2 : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 P1 : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 P0 : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 P7 : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 P6 : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 P5 : IN STD_LOGIC;
		 P4 : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 P3 : IN STD_LOGIC;
		 EQUALN : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74684_9\: COMPONENT IS true;
ATTRIBUTE noopt OF \74684_9\: COMPONENT IS true;

COMPONENT microcomputer
	PORT(n_reset : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 n_wait : IN STD_LOGIC;
		 n_int : IN STD_LOGIC;
		 n_nmi : IN STD_LOGIC;
		 n_busrq : IN STD_LOGIC;
		 dataIn : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 n_wr : OUT STD_LOGIC;
		 n_rd : OUT STD_LOGIC;
		 n_mreq : OUT STD_LOGIC;
		 n_iorq : OUT STD_LOGIC;
		 n_busak : OUT STD_LOGIC;
		 n_halt : OUT STD_LOGIC;
		 n_rfsh : OUT STD_LOGIC;
		 n_m1 : OUT STD_LOGIC;
		 address : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 dataOut : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ps2_keyboard_to_ascii
GENERIC (clk_freq : INTEGER;
			ps2_debounce_counter_size : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 ps2_clk : IN STD_LOGIC;
		 ps2_data : IN STD_LOGIC;
		 ascii_new : OUT STD_LOGIC;
		 ascii_code : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT fpga_rom
	PORT(clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT counter01_32
	PORT(clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT two_port_ram
	PORT(wren_a : IN STD_LOGIC;
		 wren_b : IN STD_LOGIC;
		 clock_a : IN STD_LOGIC;
		 clock_b : IN STD_LOGIC;
		 address_a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 address_b : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 data_a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data_b : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 q_a : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 q_b : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT spi_16bit_master
GENERIC (d_width : INTEGER;
			slaves : INTEGER
			);
	PORT(clock : IN STD_LOGIC;
		 reset_n : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 cpol : IN STD_LOGIC;
		 cpha : IN STD_LOGIC;
		 cont : IN STD_LOGIC;
		 miso : IN STD_LOGIC;
		 addr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 clk_div : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 tx_data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 sclk : OUT STD_LOGIC;
		 mosi : OUT STD_LOGIC;
		 busy : OUT STD_LOGIC;
		 rx_data : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 ss_n : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pll01_50
	PORT(inclk0 : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 c2 : OUT STD_LOGIC;
		 c3 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT fpga_rom_16k
	PORT(clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT spi_master
GENERIC (d_width : INTEGER;
			slaves : INTEGER
			);
	PORT(clock : IN STD_LOGIC;
		 reset_n : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 cpol : IN STD_LOGIC;
		 cpha : IN STD_LOGIC;
		 cont : IN STD_LOGIC;
		 miso : IN STD_LOGIC;
		 addr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 clk_div : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 tx_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 sclk : OUT STD_LOGIC;
		 mosi : OUT STD_LOGIC;
		 busy : OUT STD_LOGIC;
		 rx_data : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 ss_n : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT vga80x40
	PORT(reset : IN STD_LOGIC;
		 clk25MHz : IN STD_LOGIC;
		 FONT_D : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 ocrx : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 ocry : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 octl : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 TEXT_D : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 R : OUT STD_LOGIC;
		 G : OUT STD_LOGIC;
		 B : OUT STD_LOGIC;
		 hsync : OUT STD_LOGIC;
		 vsync : OUT STD_LOGIC;
		 cursor_x : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 cursor_y : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 FONT_A : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		 TEXT_A : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uart
GENERIC (CLOCK_DIVIDE : INTEGER;
			FLAG_HIGH : INTEGER;
			FLAG_LOW : INTEGER;
			RX_CHECK_START : INTEGER;
			RX_CHECK_STOP : INTEGER;
			RX_DELAY_RESTART : INTEGER;
			RX_ERROR : INTEGER;
			RX_IDLE : INTEGER;
			RX_READ_BITS : INTEGER;
			RX_RECEIVED : INTEGER;
			TX_DELAY_RESTART : INTEGER;
			TX_IDLE : INTEGER;
			TX_SENDING : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 rst : IN STD_LOGIC;
		 rx : IN STD_LOGIC;
		 transmit : IN STD_LOGIC;
		 data_read : IN STD_LOGIC;
		 tx_byte : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 tx : OUT STD_LOGIC;
		 received : OUT STD_LOGIC;
		 is_receiving : OUT STD_LOGIC;
		 is_transmitting : OUT STD_LOGIC;
		 recv_error : OUT STD_LOGIC;
		 data_ready : OUT STD_LOGIC;
		 rx_byte : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	10mHz :  STD_LOGIC;
SIGNAL	25Mhz :  STD_LOGIC;
SIGNAL	2mHz :  STD_LOGIC;
SIGNAL	400_KHz_CLK :  STD_LOGIC;
SIGNAL	50mHz :  STD_LOGIC;
SIGNAL	ADDRESS_LATCH :  STD_LOGIC;
SIGNAL	BAR_IN_ENABLE- :  STD_LOGIC;
SIGNAL	BOARD_INT- :  STD_LOGIC;
SIGNAL	BOARD_WAIT- :  STD_LOGIC;
SIGNAL	COUNTER_BUS :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	CPU_CLK_COUNTER :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	CTL :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CURSOR_X :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CURSOR_Y :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DATA_FROM_SDCARD :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DATA_FROM_USB_PORT :  STD_LOGIC;
SIGNAL	DATA_IN_0_A :  STD_LOGIC;
SIGNAL	DATA_IN_1_A :  STD_LOGIC;
SIGNAL	DATA_IN_2_A :  STD_LOGIC;
SIGNAL	DATA_IN_3_A :  STD_LOGIC;
SIGNAL	DATA_IN_4_A :  STD_LOGIC;
SIGNAL	DATA_IN_5_A :  STD_LOGIC;
SIGNAL	DATA_IN_6_A :  STD_LOGIC;
SIGNAL	DATA_IN_7_A :  STD_LOGIC;
SIGNAL	DATA_OUT_D0 :  STD_LOGIC;
SIGNAL	DATA_OUT_D1 :  STD_LOGIC;
SIGNAL	DATA_OUT_D2 :  STD_LOGIC;
SIGNAL	DATA_OUT_D3 :  STD_LOGIC;
SIGNAL	DATA_OUT_D4 :  STD_LOGIC;
SIGNAL	DATA_OUT_D5 :  STD_LOGIC;
SIGNAL	DATA_OUT_D6 :  STD_LOGIC;
SIGNAL	DATA_OUT_D7 :  STD_LOGIC;
SIGNAL	DATA_TO_SDCARD :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DIP_5 :  STD_LOGIC;
SIGNAL	DIP_6 :  STD_LOGIC;
SIGNAL	DIP_7 :  STD_LOGIC;
SIGNAL	DISABLE_ALL_ROM :  STD_LOGIC;
SIGNAL	END_SYNC :  STD_LOGIC;
SIGNAL	FONT_A :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	FONT_D :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	FORCE_LOW_SPEED- :  STD_LOGIC;
SIGNAL	FPGA_ROM :  STD_LOGIC;
SIGNAL	FPGA_ROM- :  STD_LOGIC;
SIGNAL	IDE_PORTA- :  STD_LOGIC;
SIGNAL	IDE_PORTB- :  STD_LOGIC;
SIGNAL	IDE_PORTC- :  STD_LOGIC;
SIGNAL	IDE_PORTCTRL- :  STD_LOGIC;
SIGNAL	IN_BOARD_RESET :  STD_LOGIC;
SIGNAL	IN_BOARD_RESET- :  STD_LOGIC;
SIGNAL	IN_CDSB- :  STD_LOGIC;
SIGNAL	IN_SDSB :  STD_LOGIC;
SIGNAL	IN_SDSB- :  STD_LOGIC;
SIGNAL	INTA_READ_DATA- :  STD_LOGIC;
SIGNAL	IO_INPUT :  STD_LOGIC;
SIGNAL	IO_OUTPUT :  STD_LOGIC;
SIGNAL	IOBYTE- :  STD_LOGIC;
SIGNAL	IOBYTE_OE- :  STD_LOGIC;
SIGNAL	JMP_ENABLE :  STD_LOGIC;
SIGNAL	JMP_ENABLE- :  STD_LOGIC;
SIGNAL	LOCAL_ADDRESS_BUS :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	LOCAL_SD_SPI_CLK :  STD_LOGIC;
SIGNAL	MEM_READ :  STD_LOGIC;
SIGNAL	MEM_WRITE :  STD_LOGIC;
SIGNAL	ocrx :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	ocry :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	OUT_CPU_CLK :  STD_LOGIC;
SIGNAL	OUT_CPU_CLK- :  STD_LOGIC;
SIGNAL	OUT_MWRT :  STD_LOGIC;
SIGNAL	OUT_pDBIN :  STD_LOGIC;
SIGNAL	OUT_pWR- :  STD_LOGIC;
SIGNAL	OUT_RAM_READ- :  STD_LOGIC;
SIGNAL	OUT_RAM_WRITE- :  STD_LOGIC;
SIGNAL	OUT_sHLTA :  STD_LOGIC;
SIGNAL	OUT_sINP :  STD_LOGIC;
SIGNAL	OUT_sINTA :  STD_LOGIC;
SIGNAL	OUT_sM1 :  STD_LOGIC;
SIGNAL	OUT_sMEMR :  STD_LOGIC;
SIGNAL	OUT_sOUT :  STD_LOGIC;
SIGNAL	OUT_sWO- :  STD_LOGIC;
SIGNAL	PORT_0- :  STD_LOGIC;
SIGNAL	PORT_1- :  STD_LOGIC;
SIGNAL	PORT_4- :  STD_LOGIC;
SIGNAL	PORT_5- :  STD_LOGIC;
SIGNAL	PORT_6- :  STD_LOGIC;
SIGNAL	PORT_7- :  STD_LOGIC;
SIGNAL	PORT_C0H- :  STD_LOGIC;
SIGNAL	PORT_C1H- :  STD_LOGIC;
SIGNAL	PORT_C2H- :  STD_LOGIC;
SIGNAL	PORT_C3H- :  STD_LOGIC;
SIGNAL	PORT_C4H- :  STD_LOGIC;
SIGNAL	PORT_C5H- :  STD_LOGIC;
SIGNAL	PORT_C6H- :  STD_LOGIC;
SIGNAL	PORT_C7H- :  STD_LOGIC;
SIGNAL	PORT_SELECT_68- :  STD_LOGIC;
SIGNAL	PORT_SELECT_69- :  STD_LOGIC;
SIGNAL	PORT_SELECT_6A- :  STD_LOGIC;
SIGNAL	PORT_SELECT_6B- :  STD_LOGIC;
SIGNAL	PORT_SELECT_6C- :  STD_LOGIC;
SIGNAL	PORT_SELECT_6D- :  STD_LOGIC;
SIGNAL	PORT_SELECT_6E- :  STD_LOGIC;
SIGNAL	PORT_SELECT_6F- :  STD_LOGIC;
SIGNAL	PRINTER_STATUS_PORT- :  STD_LOGIC;
SIGNAL	PS2_ASCII_CODE :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	PS2_DATA- :  STD_LOGIC;
SIGNAL	PS2_DATA_IN :  STD_LOGIC;
SIGNAL	PS2_KEYBOARD_STATUS :  STD_LOGIC;
SIGNAL	PS2_STATUS- :  STD_LOGIC;
SIGNAL	PS2_STATUS_IN :  STD_LOGIC;
SIGNAL	pSYNC_RAW :  STD_LOGIC;
SIGNAL	RAM_TEXT_D :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	READ_RAM :  STD_LOGIC;
SIGNAL	ROM_A12 :  STD_LOGIC;
SIGNAL	ROM_A13 :  STD_LOGIC;
SIGNAL	ROM_ADDRESS :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	ROM_OE :  STD_LOGIC;
SIGNAL	S100_A0 :  STD_LOGIC;
SIGNAL	S100_A1 :  STD_LOGIC;
SIGNAL	S100_A10 :  STD_LOGIC;
SIGNAL	S100_A11 :  STD_LOGIC;
SIGNAL	S100_A12 :  STD_LOGIC;
SIGNAL	S100_A13 :  STD_LOGIC;
SIGNAL	S100_A14 :  STD_LOGIC;
SIGNAL	S100_A15 :  STD_LOGIC;
SIGNAL	S100_A16 :  STD_LOGIC;
SIGNAL	S100_A17 :  STD_LOGIC;
SIGNAL	S100_A18 :  STD_LOGIC;
SIGNAL	S100_A19 :  STD_LOGIC;
SIGNAL	S100_A2 :  STD_LOGIC;
SIGNAL	S100_A3 :  STD_LOGIC;
SIGNAL	S100_A4 :  STD_LOGIC;
SIGNAL	S100_A5 :  STD_LOGIC;
SIGNAL	S100_A6 :  STD_LOGIC;
SIGNAL	S100_A7 :  STD_LOGIC;
SIGNAL	S100_A8 :  STD_LOGIC;
SIGNAL	S100_A9 :  STD_LOGIC;
SIGNAL	S100_INT- :  STD_LOGIC;
SIGNAL	SD_CARD_ADDRESS :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SD_CARD_BUSY :  STD_LOGIC;
SIGNAL	SD_CARD_CLK_DIV :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SD_CARD_READ_DATA- :  STD_LOGIC;
SIGNAL	SD_READ :  STD_LOGIC;
SIGNAL	SD_SLAVES :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SD_WRITE :  STD_LOGIC;
SIGNAL	SDCARD_OUT_0 :  STD_LOGIC;
SIGNAL	SDCARD_OUT_1 :  STD_LOGIC;
SIGNAL	SDCARD_OUT_2 :  STD_LOGIC;
SIGNAL	SDCARD_OUT_3 :  STD_LOGIC;
SIGNAL	SDCARD_OUT_4 :  STD_LOGIC;
SIGNAL	SDCARD_OUT_5 :  STD_LOGIC;
SIGNAL	SDCARD_OUT_6 :  STD_LOGIC;
SIGNAL	SDCARD_OUT_7 :  STD_LOGIC;
SIGNAL	SERIAL_DATA_TO_USB_PORT :  STD_LOGIC;
SIGNAL	SPI_BUSY_FLAG :  STD_LOGIC;
SIGNAL	SPI_CLK :  STD_LOGIC;
SIGNAL	SPI_CLK_DIV :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SPI_DATA_IN_BUS :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SPI_DATA_OUT_BUS :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SPI_INPUT_CS :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SPI_MASTER_CLK :  STD_LOGIC;
SIGNAL	SPI_READ :  STD_LOGIC;
SIGNAL	SPI_RTC_READ_DATA- :  STD_LOGIC;
SIGNAL	SPI_SD_CLK_SPEED :  STD_LOGIC;
SIGNAL	SPI_WRITE :  STD_LOGIC;
SIGNAL	START_BUZZER :  STD_LOGIC;
SIGNAL	START_SYNC :  STD_LOGIC;
SIGNAL	STOP_BUZZER :  STD_LOGIC;
SIGNAL	TEXT_A :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	UART_Busy :  STD_LOGIC;
SIGNAL	UART_Busy_Recieving :  STD_LOGIC;
SIGNAL	UART_Busy_Transmitting :  STD_LOGIC;
SIGNAL	UART_Byte_Recieved :  STD_LOGIC;
SIGNAL	UART_DATA_READY :  STD_LOGIC;
SIGNAL	UART_Error :  STD_LOGIC;
SIGNAL	USB_DATA- :  STD_LOGIC;
SIGNAL	USB_DATA_IN :  STD_LOGIC;
SIGNAL	USB_DATA_IN- :  STD_LOGIC;
SIGNAL	USB_DATA_IN_BUS :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	USB_DATA_OUT :  STD_LOGIC;
SIGNAL	USB_DATA_OUT_BUS :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	USB_STATUS- :  STD_LOGIC;
SIGNAL	USB_STATUS_IN :  STD_LOGIC;
SIGNAL	USB_STATUS_IN- :  STD_LOGIC;
SIGNAL	VGA_CURSOR_OE- :  STD_LOGIC;
SIGNAL	VGA_RAM_READ_DATA :  STD_LOGIC;
SIGNAL	VGA_RAM_READ_DATA- :  STD_LOGIC;
SIGNAL	VGA_RAM_SELECT :  STD_LOGIC;
SIGNAL	VGA_RAM_WRITE_DATA :  STD_LOGIC;
SIGNAL	WRITE :  STD_LOGIC;
SIGNAL	WRITE_RAM :  STD_LOGIC;
SIGNAL	Z80_ADDRESS :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	Z80_BUSAK- :  STD_LOGIC;
SIGNAL	Z80_BUSRQ- :  STD_LOGIC;
SIGNAL	Z80_HALT- :  STD_LOGIC;
SIGNAL	Z80_INTA :  STD_LOGIC;
SIGNAL	Z80_IORQ :  STD_LOGIC;
SIGNAL	Z80_IORQ- :  STD_LOGIC;
SIGNAL	Z80_LOCAL_D0 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	Z80_LOCAL_DI :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	Z80_M1 :  STD_LOGIC;
SIGNAL	Z80_M1- :  STD_LOGIC;
SIGNAL	Z80_MREQ :  STD_LOGIC;
SIGNAL	Z80_MREQ- :  STD_LOGIC;
SIGNAL	Z80_RD :  STD_LOGIC;
SIGNAL	Z80_RD- :  STD_LOGIC;
SIGNAL	Z80_RFSH- :  STD_LOGIC;
SIGNAL	Z80_WR :  STD_LOGIC;
SIGNAL	Z80_WR- :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_624 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_625 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_626 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_627 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	DFF_inst102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_628 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_629 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_630 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_631 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_632 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC_VECTOR(0 TO 7);
SIGNAL	SYNTHESIZED_WIRE_633 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_634 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_635 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_636 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_637 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC_VECTOR(0 TO 7);
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_638 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_639 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_640 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC_VECTOR(0 TO 7);
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_641 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC_VECTOR(0 TO 4);
SIGNAL	SYNTHESIZED_WIRE_642 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_643 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_644 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_645 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_646 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_647 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_648 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_649 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_650 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_651 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_652 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_653 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_654 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_655 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_168 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_656 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_171 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_173 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_657 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_658 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_659 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_660 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_661 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_662 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_663 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_664 :  STD_LOGIC_VECTOR(0 TO 1);
SIGNAL	SYNTHESIZED_WIRE_199 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_200 :  STD_LOGIC_VECTOR(0 TO 7);
SIGNAL	SYNTHESIZED_WIRE_201 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_665 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_217 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_218 :  STD_LOGIC_VECTOR(0 TO 7);
SIGNAL	SYNTHESIZED_WIRE_219 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_220 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_221 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_222 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_223 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_224 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_225 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_226 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_227 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_228 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_666 :  STD_LOGIC_VECTOR(0 TO 7);
SIGNAL	SYNTHESIZED_WIRE_667 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_668 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_669 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_238 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_239 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_670 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_240 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_242 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_243 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_244 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_245 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_246 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_671 :  STD_LOGIC_VECTOR(0 TO 6);
SIGNAL	SYNTHESIZED_WIRE_254 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_255 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_256 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_257 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_672 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_259 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_673 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_262 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_263 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_264 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_265 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_674 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_269 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_270 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_675 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_676 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_283 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_284 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_285 :  STD_LOGIC_VECTOR(0 TO 2);
SIGNAL	SYNTHESIZED_WIRE_286 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_677 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_678 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_293 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_294 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_679 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_297 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_680 :  STD_LOGIC;
SIGNAL	DFF_inst143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_305 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_306 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_307 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_309 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_311 :  STD_LOGIC;
SIGNAL	DFF_inst336 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_681 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_313 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_682 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_683 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_316 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_684 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_319 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_320 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_322 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_323 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_324 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_325 :  STD_LOGIC;
SIGNAL	DFF_inst349 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_327 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_328 :  STD_LOGIC;
SIGNAL	DFF_inst358 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_330 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_331 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_332 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_333 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_685 :  STD_LOGIC_VECTOR(0 TO 31);
SIGNAL	SYNTHESIZED_WIRE_336 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_337 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_338 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_339 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_340 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_341 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_342 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_343 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_344 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_686 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_687 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_349 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_688 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_351 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_689 :  STD_LOGIC;
SIGNAL	DFF_inst377 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_356 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_357 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_358 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_690 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_691 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_692 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_693 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_372 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_694 :  STD_LOGIC;
SIGNAL	DFF_inst387 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_377 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_378 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_379 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_695 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_381 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_696 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_697 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_698 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_699 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_700 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_701 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_702 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_703 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_422 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_426 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_427 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_704 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_445 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_705 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_706 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_462 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_464 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_465 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_466 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_467 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_468 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_469 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_470 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_707 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_472 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_476 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_478 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_479 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_480 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_481 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_482 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_483 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_484 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_708 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_486 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_709 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_710 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_711 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_712 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_713 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_714 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_497 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_715 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_500 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_503 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_505 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_506 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_716 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_511 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_717 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_513 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_718 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_719 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_535 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_720 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_721 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_722 :  STD_LOGIC;
SIGNAL	DFF_inst468 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_559 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_723 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_724 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_565 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_725 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_568 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_569 :  STD_LOGIC;
SIGNAL	DFF_inst512 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_726 :  STD_LOGIC_VECTOR(0 TO 31);
SIGNAL	SYNTHESIZED_WIRE_574 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_575 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_576 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_577 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_727 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_581 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_583 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_586 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_587 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_588 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_589 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_590 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_591 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_728 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_595 :  STD_LOGIC;
SIGNAL	DFF_inst92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_729 :  STD_LOGIC;
SIGNAL	DFF_inst97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_598 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_599 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_600 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_603 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_604 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_605 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_606 :  STD_LOGIC;
SIGNAL	DFF_inst95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_609 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_730 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_612 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_613 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_731 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_615 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_617 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_732 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_733 :  STD_LOGIC;


BEGIN 
FPGA_OUT_RAM_CS- <= '0';
FPGA_OUT_RAM_A17 <= '0';
FPGA_OUT_RAM_A18 <= '0';
LED_4 <= SD_DO;
FPGA_OUT_pHLDA <= SYNTHESIZED_WIRE_627;
PRN_ACK_LED <= DFF_inst143;
FPGA_OUT_PHANTOM <= SYNTHESIZED_WIRE_283;
P1 <= SYNTHESIZED_WIRE_535;
SD_CS_B- <= SYNTHESIZED_WIRE_719;
SD_CS_A- <= SYNTHESIZED_WIRE_716;
FPGA_OUT_IDE_RD- <= SYNTHESIZED_WIRE_171;
FPGA_OUT_IDE_WR- <= SYNTHESIZED_WIRE_173;
FPGA_OUT_8255_SEL- <= SYNTHESIZED_WIRE_656;
LED_2 <= SYNTHESIZED_WIRE_716;
LED_3 <= SYNTHESIZED_WIRE_719;
SYNTHESIZED_WIRE_1 <= '1';
SYNTHESIZED_WIRE_624 <= '1';
SYNTHESIZED_WIRE_625 <= '0';
SYNTHESIZED_WIRE_626 <= '1';
SYNTHESIZED_WIRE_19 <= '1';
SYNTHESIZED_WIRE_630 <= '0';
SYNTHESIZED_WIRE_631 <= '1';
SYNTHESIZED_WIRE_39 <= '0';
SYNTHESIZED_WIRE_44 <= '1';
SYNTHESIZED_WIRE_45 <= '0';
SYNTHESIZED_WIRE_55 <= "00000000";
SYNTHESIZED_WIRE_633 <= '0';
SYNTHESIZED_WIRE_634 <= '1';
SYNTHESIZED_WIRE_69 <= '1';
SYNTHESIZED_WIRE_636 <= '0';
SYNTHESIZED_WIRE_637 <= '1';
SYNTHESIZED_WIRE_85 <= "11111111";
SYNTHESIZED_WIRE_639 <= '0';
SYNTHESIZED_WIRE_106 <= "11111111";
SYNTHESIZED_WIRE_641 <= '0';
SYNTHESIZED_WIRE_120 <= "00000";
SYNTHESIZED_WIRE_644 <= '1';
SYNTHESIZED_WIRE_646 <= '1';
SYNTHESIZED_WIRE_142 <= '0';
SYNTHESIZED_WIRE_144 <= '0';
SYNTHESIZED_WIRE_146 <= '0';
SYNTHESIZED_WIRE_659 <= '1';
SYNTHESIZED_WIRE_661 <= '0';
SYNTHESIZED_WIRE_662 <= '1';
SYNTHESIZED_WIRE_663 <= '0';
SYNTHESIZED_WIRE_664 <= "00";
SYNTHESIZED_WIRE_200 <= "11111111";
SYNTHESIZED_WIRE_218 <= "11111111";
SYNTHESIZED_WIRE_666 <= "00000000";
SYNTHESIZED_WIRE_239 <= '1';
SYNTHESIZED_WIRE_244 <= '1';
SYNTHESIZED_WIRE_246 <= '1';
SYNTHESIZED_WIRE_671 <= "1111111";
SYNTHESIZED_WIRE_673 <= '1';
SYNTHESIZED_WIRE_674 <= '1';
SYNTHESIZED_WIRE_675 <= '0';
SYNTHESIZED_WIRE_676 <= '1';
SYNTHESIZED_WIRE_285 <= "111";
SYNTHESIZED_WIRE_294 <= '0';
SYNTHESIZED_WIRE_680 <= '1';
SYNTHESIZED_WIRE_306 <= '1';
SYNTHESIZED_WIRE_307 <= '0';
SYNTHESIZED_WIRE_682 <= '1';
SYNTHESIZED_WIRE_684 <= '1';
SYNTHESIZED_WIRE_319 <= '0';
SYNTHESIZED_WIRE_322 <= '1';
SYNTHESIZED_WIRE_323 <= '1';
SYNTHESIZED_WIRE_327 <= '1';
SYNTHESIZED_WIRE_332 <= '1';
SYNTHESIZED_WIRE_685 <= "11111111111111111111111111111111";
SYNTHESIZED_WIRE_342 <= '0';
SYNTHESIZED_WIRE_686 <= '1';
SYNTHESIZED_WIRE_349 <= '0';
SYNTHESIZED_WIRE_689 <= '1';
SYNTHESIZED_WIRE_358 <= '0';
SYNTHESIZED_WIRE_691 <= '0';
SYNTHESIZED_WIRE_692 <= '1';
SYNTHESIZED_WIRE_694 <= '1';
SYNTHESIZED_WIRE_695 <= '1';
SYNTHESIZED_WIRE_697 <= '1';
SYNTHESIZED_WIRE_700 <= '1';
SYNTHESIZED_WIRE_701 <= '0';
SYNTHESIZED_WIRE_706 <= '1';
SYNTHESIZED_WIRE_707 <= '0';
SYNTHESIZED_WIRE_709 <= '1';
SYNTHESIZED_WIRE_713 <= '1';
SYNTHESIZED_WIRE_714 <= '0';
SYNTHESIZED_WIRE_717 <= '1';
SYNTHESIZED_WIRE_720 <= '0';
SYNTHESIZED_WIRE_725 <= '1';
SYNTHESIZED_WIRE_569 <= '1';
SYNTHESIZED_WIRE_726 <= "11111111111111111111111111111111";
SYNTHESIZED_WIRE_727 <= '0';
SYNTHESIZED_WIRE_609 <= '1';
SYNTHESIZED_WIRE_730 <= '1';
SYNTHESIZED_WIRE_612 <= '1';
SYNTHESIZED_WIRE_617 <= '1';
SYNTHESIZED_WIRE_732 <= '1';



b2v_inst : microcomputer
PORT MAP(n_reset => IN_BOARD_RESET-,
		 clk => OUT_CPU_CLK,
		 n_wait => SYNTHESIZED_WIRE_0,
		 n_int => BOARD_INT-,
		 n_nmi => SYNTHESIZED_WIRE_1,
		 n_busrq => Z80_BUSRQ-,
		 dataIn => Z80_LOCAL_DI,
		 n_wr => Z80_WR-,
		 n_rd => Z80_RD-,
		 n_mreq => Z80_MREQ-,
		 n_iorq => Z80_IORQ-,
		 n_busak => Z80_BUSAK-,
		 n_halt => Z80_HALT-,
		 n_rfsh => Z80_RFSH-,
		 n_m1 => Z80_M1-,
		 address => Z80_ADDRESS,
		 dataOut => Z80_LOCAL_D0);



pSYNC_RAW <= NOT(START_SYNC OR END_SYNC OR START_SYNC OR SYNTHESIZED_WIRE_2);


FPGA_ADD_OE- <= NOT(IN_SDSB-);



FPGA_OUT_DO_OE- <= NOT(IN_SDSB-);



PROCESS(OUT_CPU_CLK,SYNTHESIZED_WIRE_624,SYNTHESIZED_WIRE_624)
BEGIN
IF (SYNTHESIZED_WIRE_624 = '0') THEN
	DFF_inst102 <= '0';
ELSIF (SYNTHESIZED_WIRE_624 = '0') THEN
	DFF_inst102 <= '1';
ELSIF (RISING_EDGE(OUT_CPU_CLK)) THEN
	DFF_inst102 <= SYNTHESIZED_WIRE_4;
END IF;
END PROCESS;


b2v_inst103 : 74165_0
PORT MAP(D => SYNTHESIZED_WIRE_625,
		 C => SYNTHESIZED_WIRE_626,
		 B => SYNTHESIZED_WIRE_626,
		 G => SYNTHESIZED_WIRE_625,
		 H => SYNTHESIZED_WIRE_625,
		 A => SYNTHESIZED_WIRE_626,
		 CLKIH => SYNTHESIZED_WIRE_625,
		 E => SYNTHESIZED_WIRE_625,
		 F => SYNTHESIZED_WIRE_625,
		 CLK => OUT_CPU_CLK-,
		 STLD => SYNTHESIZED_WIRE_15,
		 SER => SYNTHESIZED_WIRE_626,
		 QHN => SYNTHESIZED_WIRE_134);




SYNTHESIZED_WIRE_2 <= NOT(Z80_RFSH-);



FPGA_OUT_DI_OE- <= NOT(IN_SDSB-);



PROCESS(OUT_CPU_CLK-,SYNTHESIZED_WIRE_627,SYNTHESIZED_WIRE_19)
BEGIN
IF (SYNTHESIZED_WIRE_627 = '0') THEN
	SYNTHESIZED_WIRE_628 <= '0';
ELSIF (SYNTHESIZED_WIRE_19 = '0') THEN
	SYNTHESIZED_WIRE_628 <= '1';
ELSIF (RISING_EDGE(OUT_CPU_CLK-)) THEN
	SYNTHESIZED_WIRE_628 <= SYNTHESIZED_WIRE_627;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_4 <= NOT(SYNTHESIZED_WIRE_20 OR FPGA_IN_pHOLD-);



FPGA_OUT_CTL_DISABLE <= NOT(DFF_inst102);




FPGA_OUT_STATUS_DISABLE <= NOT(SYNTHESIZED_WIRE_628);



SYNTHESIZED_WIRE_627 <= NOT(Z80_BUSAK-);




b2v_inst115 : 74373_1
PORT MAP(D1 => Z80_ADDRESS(0),
		 D3 => Z80_ADDRESS(2),
		 D6 => Z80_ADDRESS(5),
		 D7 => Z80_ADDRESS(6),
		 D2 => Z80_ADDRESS(1),
		 G => ADDRESS_LATCH,
		 D4 => Z80_ADDRESS(3),
		 D5 => Z80_ADDRESS(4),
		 D8 => Z80_ADDRESS(7),
		 OEN => SYNTHESIZED_WIRE_629,
		 Q3 => S100_A2,
		 Q6 => S100_A5,
		 Q7 => S100_A6,
		 Q2 => S100_A1,
		 Q8 => S100_A7,
		 Q4 => S100_A3,
		 Q5 => S100_A4,
		 Q1 => S100_A0);


b2v_inst116 : 74373_2
PORT MAP(D1 => Z80_ADDRESS(8),
		 D3 => Z80_ADDRESS(10),
		 D6 => Z80_ADDRESS(13),
		 D7 => Z80_ADDRESS(14),
		 D2 => Z80_ADDRESS(9),
		 G => ADDRESS_LATCH,
		 D4 => Z80_ADDRESS(11),
		 D5 => Z80_ADDRESS(12),
		 D8 => Z80_ADDRESS(15),
		 OEN => SYNTHESIZED_WIRE_629,
		 Q3 => SYNTHESIZED_WIRE_581,
		 Q6 => SYNTHESIZED_WIRE_102,
		 Q7 => SYNTHESIZED_WIRE_100,
		 Q2 => SYNTHESIZED_WIRE_583,
		 Q8 => SYNTHESIZED_WIRE_105,
		 Q4 => SYNTHESIZED_WIRE_586,
		 Q5 => SYNTHESIZED_WIRE_96,
		 Q1 => SYNTHESIZED_WIRE_577);


b2v_inst117 : 74373_3
PORT MAP(D1 => SYNTHESIZED_WIRE_630,
		 D3 => SYNTHESIZED_WIRE_630,
		 D6 => SYNTHESIZED_WIRE_630,
		 D7 => SYNTHESIZED_WIRE_630,
		 D2 => SYNTHESIZED_WIRE_630,
		 G => ADDRESS_LATCH,
		 D4 => SYNTHESIZED_WIRE_630,
		 D5 => SYNTHESIZED_WIRE_630,
		 D8 => SYNTHESIZED_WIRE_630,
		 OEN => SYNTHESIZED_WIRE_629,
		 Q3 => S100_A18,
		 Q2 => S100_A17,
		 Q4 => S100_A19,
		 Q1 => S100_A16);


SYNTHESIZED_WIRE_615 <= NOT(SYNTHESIZED_WIRE_32);





SYNTHESIZED_WIRE_15 <= NOT(pSYNC_RAW AND Z80_IORQ);


b2v_inst121 : 74165_4
PORT MAP(D => SYNTHESIZED_WIRE_631,
		 C => SYNTHESIZED_WIRE_631,
		 B => SYNTHESIZED_WIRE_631,
		 G => SYNTHESIZED_WIRE_631,
		 H => SYNTHESIZED_WIRE_631,
		 A => SYNTHESIZED_WIRE_631,
		 CLKIH => SYNTHESIZED_WIRE_39,
		 E => SYNTHESIZED_WIRE_631,
		 F => SYNTHESIZED_WIRE_631,
		 CLK => OUT_CPU_CLK-,
		 STLD => SYNTHESIZED_WIRE_42,
		 SER => SYNTHESIZED_WIRE_631,
		 QHN => SYNTHESIZED_WIRE_645);




PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_44,SYNTHESIZED_WIRE_46)
BEGIN
IF (SYNTHESIZED_WIRE_44 = '0') THEN
	JMP_ENABLE- <= '0';
ELSIF (SYNTHESIZED_WIRE_46 = '0') THEN
	JMP_ENABLE- <= '1';
ELSIF (RISING_EDGE(IN_BOARD_RESET-)) THEN
	JMP_ENABLE- <= SYNTHESIZED_WIRE_45;
END IF;
END PROCESS;


PROCESS(FPGA_IN_DI0,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(0) <= FPGA_IN_DI0;
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_IN_DI1,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(1) <= FPGA_IN_DI1;
ELSE
	Z80_LOCAL_DI(1) <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_IN_DI2,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(2) <= FPGA_IN_DI2;
ELSE
	Z80_LOCAL_DI(2) <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_IN_DI3,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(3) <= FPGA_IN_DI3;
ELSE
	Z80_LOCAL_DI(3) <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_IN_DI4,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(4) <= FPGA_IN_DI4;
ELSE
	Z80_LOCAL_DI(4) <= 'Z';
END IF;
END PROCESS;


ADDRESS_LATCH <= NOT(pSYNC_RAW AND OUT_CPU_CLK-);


PROCESS(FPGA_IN_DI5,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(5) <= FPGA_IN_DI5;
ELSE
	Z80_LOCAL_DI(5) <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_IN_DI6,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(6) <= FPGA_IN_DI6;
ELSE
	Z80_LOCAL_DI(6) <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_IN_DI7,SYNTHESIZED_WIRE_632)
BEGIN
if (SYNTHESIZED_WIRE_632 = '1') THEN
	Z80_LOCAL_DI(7) <= FPGA_IN_DI7;
ELSE
	Z80_LOCAL_DI(7) <= 'Z';
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(7) <= SYNTHESIZED_WIRE_55(0);
ELSE
	Z80_LOCAL_DI(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(6) <= SYNTHESIZED_WIRE_55(1);
ELSE
	Z80_LOCAL_DI(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(5) <= SYNTHESIZED_WIRE_55(2);
ELSE
	Z80_LOCAL_DI(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(4) <= SYNTHESIZED_WIRE_55(3);
ELSE
	Z80_LOCAL_DI(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(3) <= SYNTHESIZED_WIRE_55(4);
ELSE
	Z80_LOCAL_DI(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(2) <= SYNTHESIZED_WIRE_55(5);
ELSE
	Z80_LOCAL_DI(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(1) <= SYNTHESIZED_WIRE_55(6);
ELSE
	Z80_LOCAL_DI(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_55,JMP_ENABLE)
BEGIN
if (JMP_ENABLE = '1') THEN
	Z80_LOCAL_DI(0) <= SYNTHESIZED_WIRE_55(7);
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(DATA_OUT_D2,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D2 <= DATA_OUT_D2;
ELSE
	FPGA_BI_D2 <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_BI_D2,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(2) <= FPGA_BI_D2;
ELSE
	Z80_LOCAL_DI(2) <= 'Z';
END IF;
END PROCESS;


PROCESS(DATA_OUT_D3,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D3 <= DATA_OUT_D3;
ELSE
	FPGA_BI_D3 <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_BI_D3,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(3) <= FPGA_BI_D3;
ELSE
	Z80_LOCAL_DI(3) <= 'Z';
END IF;
END PROCESS;


b2v_inst138 : 74684_5
PORT MAP(P2 => SYNTHESIZED_WIRE_633,
		 Q2 => SYNTHESIZED_WIRE_633,
		 P1 => SYNTHESIZED_WIRE_633,
		 Q1 => SYNTHESIZED_WIRE_633,
		 P0 => SYNTHESIZED_WIRE_633,
		 Q0 => SYNTHESIZED_WIRE_633,
		 P7 => S100_A7,
		 Q7 => SYNTHESIZED_WIRE_633,
		 Q6 => SYNTHESIZED_WIRE_633,
		 P6 => S100_A6,
		 Q5 => SYNTHESIZED_WIRE_634,
		 P5 => S100_A5,
		 P4 => S100_A4,
		 Q4 => SYNTHESIZED_WIRE_634,
		 Q3 => SYNTHESIZED_WIRE_633,
		 P3 => S100_A3,
		 EQUALN => SYNTHESIZED_WIRE_638);



FPGA_OUT_HIGH_ROM_LED- <= SYNTHESIZED_WIRE_67 OR DISABLE_ALL_ROM;


PROCESS(DATA_OUT_D4,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D4 <= DATA_OUT_D4;
ELSE
	FPGA_BI_D4 <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_BI_D4,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(4) <= FPGA_BI_D4;
ELSE
	Z80_LOCAL_DI(4) <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_669 <= PORT_C1H- OR SYNTHESIZED_WIRE_635;


PROCESS(IN_BOARD_RESET-,FPGA_IN_PRN_ACK,SYNTHESIZED_WIRE_70)
BEGIN
IF (FPGA_IN_PRN_ACK = '0') THEN
	DFF_inst143 <= '0';
ELSIF (SYNTHESIZED_WIRE_70 = '0') THEN
	DFF_inst143 <= '1';
ELSIF (RISING_EDGE(IN_BOARD_RESET-)) THEN
	DFF_inst143 <= SYNTHESIZED_WIRE_69;
END IF;
END PROCESS;



PROCESS(DATA_OUT_D5,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D5 <= DATA_OUT_D5;
ELSE
	FPGA_BI_D5 <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_BI_D5,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(5) <= FPGA_BI_D5;
ELSE
	Z80_LOCAL_DI(5) <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_238 <= NOT(IOBYTE- OR SYNTHESIZED_WIRE_71);


SYNTHESIZED_WIRE_283 <= VGA_RAM_WRITE_DATA OR VGA_RAM_READ_DATA;


b2v_inst149 : 74684_6
PORT MAP(P2 => SYNTHESIZED_WIRE_636,
		 Q2 => SYNTHESIZED_WIRE_636,
		 P1 => SYNTHESIZED_WIRE_636,
		 Q1 => SYNTHESIZED_WIRE_636,
		 P0 => SYNTHESIZED_WIRE_636,
		 Q0 => SYNTHESIZED_WIRE_636,
		 P7 => S100_A15,
		 Q7 => SYNTHESIZED_WIRE_637,
		 Q6 => SYNTHESIZED_WIRE_637,
		 P6 => S100_A14,
		 Q5 => SYNTHESIZED_WIRE_637,
		 P5 => S100_A13,
		 P4 => S100_A12,
		 Q4 => SYNTHESIZED_WIRE_637,
		 Q3 => SYNTHESIZED_WIRE_636,
		 P3 => SYNTHESIZED_WIRE_636,
		 EQUALN => SYNTHESIZED_WIRE_665);


USB_TX_BUSY_LED <= NOT(UART_Busy);



PROCESS(DATA_OUT_D6,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D6 <= DATA_OUT_D6;
ELSE
	FPGA_BI_D6 <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_BI_D6,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(6) <= FPGA_BI_D6;
ELSE
	Z80_LOCAL_DI(6) <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_84 <= NOT(UART_Busy_Transmitting);



SYNTHESIZED_WIRE_331 <= SYNTHESIZED_WIRE_84 AND IN_BOARD_RESET-;



PROCESS(DATA_OUT_D7,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D7 <= DATA_OUT_D7;
ELSE
	FPGA_BI_D7 <= 'Z';
END IF;
END PROCESS;


PROCESS(FPGA_BI_D7,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(7) <= FPGA_BI_D7;
ELSE
	Z80_LOCAL_DI(7) <= 'Z';
END IF;
END PROCESS;



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_85,USB_DATA_OUT,Z80_LOCAL_D0)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	USB_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_85 = '0') THEN
	USB_DATA_OUT_BUS <= '1';
ELSIF (USB_DATA_OUT = '1') THEN
	USB_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(7) <= SYNTHESIZED_WIRE_86(7);
ELSE
	Z80_LOCAL_DI(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(6) <= SYNTHESIZED_WIRE_86(6);
ELSE
	Z80_LOCAL_DI(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(5) <= SYNTHESIZED_WIRE_86(5);
ELSE
	Z80_LOCAL_DI(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(4) <= SYNTHESIZED_WIRE_86(4);
ELSE
	Z80_LOCAL_DI(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(3) <= SYNTHESIZED_WIRE_86(3);
ELSE
	Z80_LOCAL_DI(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(2) <= SYNTHESIZED_WIRE_86(2);
ELSE
	Z80_LOCAL_DI(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(1) <= SYNTHESIZED_WIRE_86(1);
ELSE
	Z80_LOCAL_DI(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_86,USB_DATA_IN)
BEGIN
if (USB_DATA_IN = '1') THEN
	Z80_LOCAL_DI(0) <= SYNTHESIZED_WIRE_86(0);
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;


b2v_inst16 : 74138_7
PORT MAP(A => S100_A0,
		 B => S100_A1,
		 G1 => SYNTHESIZED_WIRE_87,
		 C => S100_A2,
		 G2AN => SYNTHESIZED_WIRE_638,
		 G2BN => SYNTHESIZED_WIRE_638,
		 Y0N => IDE_PORTA-,
		 Y1N => IDE_PORTB-,
		 Y2N => IDE_PORTC-,
		 Y3N => IDE_PORTCTRL-,
		 Y4N => USB_STATUS-,
		 Y5N => USB_DATA-,
		 Y6N => IOBYTE-);


SYNTHESIZED_WIRE_264 <= IN_BOARD_RESET- AND PS2_DATA-;



b2v_inst162 : ps2_keyboard_to_ascii
GENERIC MAP(clk_freq => 50000000,
			ps2_debounce_counter_size => 8
			)
PORT MAP(clk => 50mHz,
		 ps2_clk => FPGA_IN_PS2_CLK,
		 ps2_data => FPGA_IN_PS2_DATA,
		 ascii_new => SYNTHESIZED_WIRE_265,
		 ascii_code => PS2_ASCII_CODE);


SYNTHESIZED_WIRE_632 <= SYNTHESIZED_WIRE_90 AND SYNTHESIZED_WIRE_91 AND SYNTHESIZED_WIRE_92 AND IOBYTE_OE- AND OUT_pDBIN AND OUT_sINP AND SYNTHESIZED_WIRE_93 AND SYNTHESIZED_WIRE_94;


USB_DATA_OUT <= NOT(USB_DATA- OR OUT_pWR-);


SYNTHESIZED_WIRE_305 <= NOT(SYNTHESIZED_WIRE_95 OR OUT_pWR- OR PORT_7-);


SYNTHESIZED_WIRE_657 <= FPGA_IN_PRN_ACK AND IN_BOARD_RESET-;


SYNTHESIZED_WIRE_257 <= DIP_7 AND FORCE_LOW_SPEED-;


b2v_inst168 : 74157_8
PORT MAP(A1 => SYNTHESIZED_WIRE_96,
		 B1 => SYNTHESIZED_WIRE_639,
		 SEL => SYNTHESIZED_WIRE_640,
		 B2 => SYNTHESIZED_WIRE_639,
		 A3 => SYNTHESIZED_WIRE_100,
		 B3 => SYNTHESIZED_WIRE_639,
		 A2 => SYNTHESIZED_WIRE_102,
		 B4 => SYNTHESIZED_WIRE_639,
		 GN => SYNTHESIZED_WIRE_639,
		 A4 => SYNTHESIZED_WIRE_105,
		 Y2 => S100_A13,
		 Y1 => S100_A12,
		 Y4 => S100_A15,
		 Y3 => S100_A14);



SYNTHESIZED_WIRE_642 <= NOT(OUT_pDBIN);



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_106,USB_DATA_IN,USB_DATA_IN_BUS)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_86 <= '0';
ELSIF (SYNTHESIZED_WIRE_106 = '0') THEN
	SYNTHESIZED_WIRE_86 <= '1';
ELSIF (USB_DATA_IN = '1') THEN
	SYNTHESIZED_WIRE_86 <= USB_DATA_IN_BUS;
END IF;
END PROCESS;



PROCESS(SYNTHESIZED_WIRE_107,PS2_STATUS_IN)
BEGIN
if (PS2_STATUS_IN = '1') THEN
	Z80_LOCAL_DI(0) <= SYNTHESIZED_WIRE_107;
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_108,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(6) <= SYNTHESIZED_WIRE_108(6);
ELSE
	Z80_LOCAL_DI(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_108,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(5) <= SYNTHESIZED_WIRE_108(5);
ELSE
	Z80_LOCAL_DI(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_108,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(4) <= SYNTHESIZED_WIRE_108(4);
ELSE
	Z80_LOCAL_DI(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_108,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(3) <= SYNTHESIZED_WIRE_108(3);
ELSE
	Z80_LOCAL_DI(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_108,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(2) <= SYNTHESIZED_WIRE_108(2);
ELSE
	Z80_LOCAL_DI(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_108,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(1) <= SYNTHESIZED_WIRE_108(1);
ELSE
	Z80_LOCAL_DI(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_108,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(0) <= SYNTHESIZED_WIRE_108(0);
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;



SYNTHESIZED_WIRE_160 <= OUT_sINP OR OUT_sOUT;


b2v_inst176 : 74684_9
PORT MAP(P2 => SYNTHESIZED_WIRE_641,
		 Q2 => SYNTHESIZED_WIRE_641,
		 P1 => SYNTHESIZED_WIRE_641,
		 Q1 => SYNTHESIZED_WIRE_641,
		 P0 => SYNTHESIZED_WIRE_641,
		 Q0 => SYNTHESIZED_WIRE_641,
		 P7 => S100_A7,
		 Q7 => SYNTHESIZED_WIRE_641,
		 Q6 => SYNTHESIZED_WIRE_641,
		 P6 => S100_A6,
		 Q5 => SYNTHESIZED_WIRE_641,
		 P5 => S100_A5,
		 P4 => S100_A4,
		 Q4 => SYNTHESIZED_WIRE_641,
		 Q3 => SYNTHESIZED_WIRE_641,
		 P3 => S100_A3,
		 EQUALN => SYNTHESIZED_WIRE_651);


SYNTHESIZED_WIRE_629 <= NOT(IN_SDSB-);



SYNTHESIZED_WIRE_591 <= NOT(IN_SDSB-);



CTL(7 DOWNTO 3) <= NOT(SYNTHESIZED_WIRE_120);



b2v_inst18 : 74373_10
PORT MAP(D1 => DIP7,
		 D3 => DIP5,
		 D6 => DIP_5,
		 D7 => DIP_6,
		 D2 => DIP6,
		 G => SYNTHESIZED_WIRE_642,
		 D4 => DIP4,
		 D5 => DIP3,
		 D8 => DIP_7,
		 OEN => IOBYTE_OE-,
		 Q3 => Z80_LOCAL_DI(2),
		 Q6 => Z80_LOCAL_DI(5),
		 Q7 => Z80_LOCAL_DI(6),
		 Q2 => Z80_LOCAL_DI(1),
		 Q8 => Z80_LOCAL_DI(7),
		 Q4 => Z80_LOCAL_DI(3),
		 Q5 => Z80_LOCAL_DI(4),
		 Q1 => Z80_LOCAL_DI(0));




PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_647 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_647 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_647 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(1))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_648 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_648 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_648 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(2))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_649 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_649 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_649 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(3))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_650 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_650 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_650 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(4))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_652 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_652 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_652 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_163 <= NOT(OUT_sOUT);



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(5))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_654 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_654 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_654 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_137 <= NOT(OUT_pDBIN);



BOARD_WAIT- <= NOT(SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_645 OR SYNTHESIZED_WIRE_645);


USB_DATA_IN <= NOT(USB_DATA- OR SYNTHESIZED_WIRE_137);


SYNTHESIZED_WIRE_149 <= NOT(OUT_pDBIN);




UART_Busy <= UART_Busy_Transmitting OR UART_Busy_Transmitting;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,UART_DATA_READY)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_221 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_221 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_221 <= UART_DATA_READY;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,UART_Busy)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_219 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_219 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_219 <= UART_Busy;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,UART_Byte_Recieved)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_222 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_222 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_222 <= UART_Byte_Recieved;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,UART_Busy_Recieving)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_220 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_220 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_220 <= UART_Busy_Recieving;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,SYNTHESIZED_WIRE_142)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_224 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_224 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_224 <= SYNTHESIZED_WIRE_142;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,SYNTHESIZED_WIRE_144)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_226 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_226 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_226 <= SYNTHESIZED_WIRE_144;
END IF;
END PROCESS;


WRITE_RAM <= NOT(JMP_ENABLE OR OUT_RAM_WRITE-);



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,SYNTHESIZED_WIRE_146)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_223 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_223 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_223 <= SYNTHESIZED_WIRE_146;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_646,USB_STATUS_IN,UART_Error)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_225 <= '0';
ELSIF (SYNTHESIZED_WIRE_646 = '0') THEN
	SYNTHESIZED_WIRE_225 <= '1';
ELSIF (USB_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_225 <= UART_Error;
END IF;
END PROCESS;




SYNTHESIZED_WIRE_87 <= OUT_sINP OR OUT_sOUT;


USB_STATUS_IN <= NOT(USB_STATUS- OR SYNTHESIZED_WIRE_149);


USB_STATUS_IN- <= NOT(USB_STATUS_IN);



SYNTHESIZED_WIRE_513 <= OUT_sINP OR OUT_sOUT;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(6))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_653 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_653 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_653 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_644,SYNTHESIZED_WIRE_643,Z80_LOCAL_D0(7))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_655 <= '0';
ELSIF (SYNTHESIZED_WIRE_644 = '0') THEN
	SYNTHESIZED_WIRE_655 <= '1';
ELSIF (SYNTHESIZED_WIRE_643 = '1') THEN
	SYNTHESIZED_WIRE_655 <= Z80_LOCAL_D0;
END IF;
END PROCESS;



PROCESS(SYNTHESIZED_WIRE_154,PS2_DATA_IN)
BEGIN
if (PS2_DATA_IN = '1') THEN
	Z80_LOCAL_DI(7) <= SYNTHESIZED_WIRE_154;
ELSE
	Z80_LOCAL_DI(7) <= 'Z';
END IF;
END PROCESS;



F_BAR0 <= NOT(SYNTHESIZED_WIRE_647);



PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(7) <= SYNTHESIZED_WIRE_156(7);
ELSE
	Z80_LOCAL_DI(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(6) <= SYNTHESIZED_WIRE_156(6);
ELSE
	Z80_LOCAL_DI(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(5) <= SYNTHESIZED_WIRE_156(5);
ELSE
	Z80_LOCAL_DI(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(4) <= SYNTHESIZED_WIRE_156(4);
ELSE
	Z80_LOCAL_DI(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(3) <= SYNTHESIZED_WIRE_156(3);
ELSE
	Z80_LOCAL_DI(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(2) <= SYNTHESIZED_WIRE_156(2);
ELSE
	Z80_LOCAL_DI(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(1) <= SYNTHESIZED_WIRE_156(1);
ELSE
	Z80_LOCAL_DI(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_156,VGA_RAM_READ_DATA)
BEGIN
if (VGA_RAM_READ_DATA = '1') THEN
	Z80_LOCAL_DI(0) <= SYNTHESIZED_WIRE_156(0);
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;


F_BAR1 <= NOT(SYNTHESIZED_WIRE_648);



F_BAR2 <= NOT(SYNTHESIZED_WIRE_649);



F_BAR3 <= NOT(SYNTHESIZED_WIRE_650);



b2v_inst217 : 74138_11
PORT MAP(A => S100_A0,
		 B => S100_A1,
		 G1 => SYNTHESIZED_WIRE_160,
		 C => S100_A2,
		 G2AN => SYNTHESIZED_WIRE_651,
		 G2BN => SYNTHESIZED_WIRE_651,
		 Y0N => PORT_0-,
		 Y2N => PS2_STATUS-,
		 Y3N => PS2_DATA-,
		 Y6N => PORT_6-,
		 Y7N => PORT_7-);


SYNTHESIZED_WIRE_643 <= NOT(OUT_pWR- OR SYNTHESIZED_WIRE_163 OR PORT_6-);


F_BAR4 <= NOT(SYNTHESIZED_WIRE_652);



USB_RX_BUSY_LED <= NOT(UART_Byte_Recieved);



F_BAR6 <= NOT(SYNTHESIZED_WIRE_653);



F_BAR5 <= NOT(SYNTHESIZED_WIRE_654);



F_BAR7 <= NOT(SYNTHESIZED_WIRE_655);



SYNTHESIZED_WIRE_46 <= NOT(MEM_READ AND SYNTHESIZED_WIRE_168);


SYNTHESIZED_WIRE_173 <= NOT(SYNTHESIZED_WIRE_169 AND OUT_sOUT);


SYNTHESIZED_WIRE_171 <= NOT(OUT_sINP AND OUT_pDBIN);


SYNTHESIZED_WIRE_169 <= NOT(OUT_pWR-);



SYNTHESIZED_WIRE_656 <= IDE_PORTA- AND IDE_PORTB- AND IDE_PORTC- AND IDE_PORTCTRL-;


5V_OUT_IDE_PORTS_RD- <= SYNTHESIZED_WIRE_656 OR SYNTHESIZED_WIRE_171;


5V_OUT_IDE_PORTS_WR- <= SYNTHESIZED_WIRE_656 OR SYNTHESIZED_WIRE_173;


DATA_OUT_D0 <= Z80_LOCAL_D0(0) OR Z80_LOCAL_D0(0);



PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(0))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_0 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_0 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_0 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_678 <= PORT_C2H- OR SYNTHESIZED_WIRE_660;


PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(1))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_1 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_1 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_1 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(2))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_2 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_2 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_2 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


b2v_inst235 : 74684_12
PORT MAP(P2 => SYNTHESIZED_WIRE_661,
		 Q2 => SYNTHESIZED_WIRE_661,
		 P1 => SYNTHESIZED_WIRE_661,
		 Q1 => SYNTHESIZED_WIRE_661,
		 P0 => SYNTHESIZED_WIRE_661,
		 Q0 => SYNTHESIZED_WIRE_661,
		 P7 => S100_A7,
		 Q7 => SYNTHESIZED_WIRE_662,
		 Q6 => SYNTHESIZED_WIRE_662,
		 P6 => S100_A6,
		 Q5 => SYNTHESIZED_WIRE_661,
		 P5 => S100_A5,
		 P4 => S100_A4,
		 Q4 => SYNTHESIZED_WIRE_661,
		 Q3 => SYNTHESIZED_WIRE_661,
		 P3 => S100_A3,
		 EQUALN => SYNTHESIZED_WIRE_718);


SYNTHESIZED_WIRE_635 <= NOT(OUT_pDBIN);



CURSOR_X(7) <= SYNTHESIZED_WIRE_663 OR SYNTHESIZED_WIRE_663;


CURSOR_Y(7 DOWNTO 6) <= SYNTHESIZED_WIRE_664 OR SYNTHESIZED_WIRE_664;



DATA_OUT_D1 <= Z80_LOCAL_D0(1) OR Z80_LOCAL_D0(1);


b2v_inst240 : fpga_rom
PORT MAP(clock => 25Mhz,
		 address => FONT_A,
		 q => FONT_D);


IN_BOARD_RESET <= NOT(IN_BOARD_RESET-);




PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_200,SYNTHESIZED_WIRE_199,Z80_LOCAL_D0)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	ocrx <= '0';
ELSIF (SYNTHESIZED_WIRE_200 = '0') THEN
	ocrx <= '1';
ELSIF (SYNTHESIZED_WIRE_199 = '1') THEN
	ocrx <= Z80_LOCAL_D0;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_201 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_199 <= NOT(OUT_pWR- OR SYNTHESIZED_WIRE_201 OR PORT_C0H-);



SYNTHESIZED_WIRE_168 <= NOT(SYNTHESIZED_WIRE_665);



PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(3))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_3 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_3 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_3 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


DATA_OUT_D2 <= Z80_LOCAL_D0(2) OR Z80_LOCAL_D0(2);


b2v_inst250 : counter01_32
PORT MAP(clock => OUT_CPU_CLK,
		 q => CPU_CLK_COUNTER);


PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(4))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_4 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_4 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_4 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


b2v_inst252 : 74244_13
PORT MAP(1A2 => SYNTHESIZED_WIRE_648,
		 1A4 => SYNTHESIZED_WIRE_650,
		 1A1 => SYNTHESIZED_WIRE_647,
		 1A3 => SYNTHESIZED_WIRE_649,
		 1GN => BAR_IN_ENABLE-,
		 2A3 => SYNTHESIZED_WIRE_653,
		 2GN => BAR_IN_ENABLE-,
		 2A1 => SYNTHESIZED_WIRE_652,
		 2A4 => SYNTHESIZED_WIRE_655,
		 2A2 => SYNTHESIZED_WIRE_654,
		 1Y2 => Z80_LOCAL_DI(1),
		 1Y4 => Z80_LOCAL_DI(3),
		 2Y1 => Z80_LOCAL_DI(4),
		 1Y1 => Z80_LOCAL_DI(0),
		 2Y3 => Z80_LOCAL_DI(6),
		 2Y4 => Z80_LOCAL_DI(7),
		 1Y3 => Z80_LOCAL_DI(2),
		 2Y2 => Z80_LOCAL_DI(5));


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_218,SYNTHESIZED_WIRE_217,Z80_LOCAL_D0)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	ocry <= '0';
ELSIF (SYNTHESIZED_WIRE_218 = '0') THEN
	ocry <= '1';
ELSIF (SYNTHESIZED_WIRE_217 = '1') THEN
	ocry <= Z80_LOCAL_D0;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_227 <= NOT(PORT_6-);



b2v_inst255 : 74244_14
PORT MAP(1A2 => SYNTHESIZED_WIRE_219,
		 1A4 => SYNTHESIZED_WIRE_220,
		 1A1 => SYNTHESIZED_WIRE_221,
		 1A3 => SYNTHESIZED_WIRE_222,
		 1GN => USB_STATUS_IN-,
		 2A3 => SYNTHESIZED_WIRE_223,
		 2GN => USB_STATUS_IN-,
		 2A1 => SYNTHESIZED_WIRE_224,
		 2A4 => SYNTHESIZED_WIRE_225,
		 2A2 => SYNTHESIZED_WIRE_226,
		 1Y2 => Z80_LOCAL_DI(1),
		 1Y4 => Z80_LOCAL_DI(3),
		 2Y1 => Z80_LOCAL_DI(4),
		 1Y1 => Z80_LOCAL_DI(0),
		 2Y3 => Z80_LOCAL_DI(6),
		 2Y4 => Z80_LOCAL_DI(7),
		 1Y3 => Z80_LOCAL_DI(2),
		 2Y2 => Z80_LOCAL_DI(5));


BAR_IN_ENABLE- <= NOT(OUT_pDBIN AND OUT_sINP AND SYNTHESIZED_WIRE_227);


SYNTHESIZED_WIRE_228 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_217 <= NOT(OUT_pWR- OR SYNTHESIZED_WIRE_228 OR PORT_C1H-);


SYNTHESIZED_WIRE_242 <= SYNTHESIZED_WIRE_666 OR SYNTHESIZED_WIRE_666;


DATA_OUT_D3 <= Z80_LOCAL_D0(3) OR Z80_LOCAL_D0(3);


b2v_inst260 : 74373b_15
PORT MAP(G => SYNTHESIZED_WIRE_667,
		 OEN => SYNTHESIZED_WIRE_668,
		 D => CURSOR_X,
		 Q => Z80_LOCAL_DI);


b2v_inst261 : 74373b_16
PORT MAP(G => SYNTHESIZED_WIRE_635,
		 OEN => SYNTHESIZED_WIRE_669,
		 D => CURSOR_Y,
		 Q => Z80_LOCAL_DI);


PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(5))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_5 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_5 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_5 <= Z80_LOCAL_D0;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_640 <= OUT_sINP OR OUT_sOUT;



PROCESS(SYNTHESIZED_WIRE_238,IN_BOARD_RESET-,SYNTHESIZED_WIRE_239)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_670 <= '0';
ELSIF (SYNTHESIZED_WIRE_239 = '0') THEN
	SYNTHESIZED_WIRE_670 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_238)) THEN
	SYNTHESIZED_WIRE_670 <= Z80_LOCAL_D0(0);
END IF;
END PROCESS;


SYNTHESIZED_WIRE_240 <= NOT(S100_A15);



FPGA_OUT_RAM_A16 <= SYNTHESIZED_WIRE_670 AND SYNTHESIZED_WIRE_240;



DATA_OUT_D4 <= Z80_LOCAL_D0(4) OR Z80_LOCAL_D0(4);


FPGA_OUT_HIGH_RAM_LED- <= NOT(SYNTHESIZED_WIRE_670);



b2v_inst271 : two_port_ram
PORT MAP(wren_a => VGA_RAM_WRITE_DATA,
		 wren_b => SYNTHESIZED_WIRE_666,
		 clock_a => 25Mhz,
		 clock_b => 25Mhz,
		 address_a => LOCAL_ADDRESS_BUS(11 DOWNTO 0),
		 address_b => TEXT_A,
		 data_a => Z80_LOCAL_D0,
		 data_b => SYNTHESIZED_WIRE_242,
		 q_a => SYNTHESIZED_WIRE_156,
		 q_b => RAM_TEXT_D);


PROCESS(SYNTHESIZED_WIRE_243,IN_BOARD_RESET-,SYNTHESIZED_WIRE_244)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DISABLE_ALL_ROM <= '0';
ELSIF (SYNTHESIZED_WIRE_244 = '0') THEN
	DISABLE_ALL_ROM <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_243)) THEN
	DISABLE_ALL_ROM <= Z80_LOCAL_D0(1);
END IF;
END PROCESS;


SYNTHESIZED_WIRE_445 <= NOT(OUT_sOUT);



PROCESS(SYNTHESIZED_WIRE_245,IN_BOARD_RESET-,SYNTHESIZED_WIRE_246)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	ROM_A12 <= '0';
ELSIF (SYNTHESIZED_WIRE_246 = '0') THEN
	ROM_A12 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_245)) THEN
	ROM_A12 <= Z80_LOCAL_D0(0);
END IF;
END PROCESS;



PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(6))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_6 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_6 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_6 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_671,PS2_DATA_IN,PS2_ASCII_CODE)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_108 <= '0';
ELSIF (SYNTHESIZED_WIRE_671 = '0') THEN
	SYNTHESIZED_WIRE_108 <= '1';
ELSIF (PS2_DATA_IN = '1') THEN
	SYNTHESIZED_WIRE_108 <= PS2_ASCII_CODE;
END IF;
END PROCESS;



PROCESS(SYNTHESIZED_WIRE_657,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_658,Z80_LOCAL_D0(7))
BEGIN
IF (SYNTHESIZED_WIRE_657 = '0') THEN
	FPGA_OUT_PRN_7 <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_7 <= '1';
ELSIF (SYNTHESIZED_WIRE_658 = '1') THEN
	FPGA_OUT_PRN_7 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


DATA_OUT_D5 <= Z80_LOCAL_D0(5) OR Z80_LOCAL_D0(5);


b2v_inst280 : 74373b_17
PORT MAP(G => ADDRESS_LATCH,
		 OEN => SYNTHESIZED_WIRE_254,
		 D => Z80_ADDRESS(7 DOWNTO 0),
		 Q => LOCAL_ADDRESS_BUS(7 DOWNTO 0));


SYNTHESIZED_WIRE_254 <= NOT(IN_SDSB-);



b2v_inst282 : 74373b_18
PORT MAP(G => ADDRESS_LATCH,
		 OEN => SYNTHESIZED_WIRE_255,
		 D => Z80_ADDRESS(15 DOWNTO 8),
		 Q => LOCAL_ADDRESS_BUS(15 DOWNTO 8));


SYNTHESIZED_WIRE_255 <= NOT(IN_SDSB-);



SYNTHESIZED_WIRE_259 <= NOT(OUT_MWRT AND VGA_RAM_SELECT);


SYNTHESIZED_WIRE_42 <= NOT(Z80_MREQ AND SYNTHESIZED_WIRE_256 AND pSYNC_RAW);


SYNTHESIZED_WIRE_256 <= NOT(FPGA_ROM-);



b2v_inst287 : 21mux_19
PORT MAP(S => SYNTHESIZED_WIRE_257,
		 B => 2mHz,
		 A => 25Mhz,
		 Y => OUT_CPU_CLK);


SYNTHESIZED_WIRE_427 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_71 <= NOT(IO_OUTPUT);



SYNTHESIZED_WIRE_731 <= NOT(Z80_RD- AND SYNTHESIZED_WIRE_672);


VGA_RAM_WRITE_DATA <= NOT(SYNTHESIZED_WIRE_259 OR OUT_pWR-);


SYNTHESIZED_WIRE_20 <= NOT(SYNTHESIZED_WIRE_628);



PROCESS(OUT_CPU_CLK,SYNTHESIZED_WIRE_673,SYNTHESIZED_WIRE_673)
BEGIN
IF (SYNTHESIZED_WIRE_673 = '0') THEN
	Z80_BUSRQ- <= '0';
ELSIF (SYNTHESIZED_WIRE_673 = '0') THEN
	Z80_BUSRQ- <= '1';
ELSIF (RISING_EDGE(OUT_CPU_CLK)) THEN
	Z80_BUSRQ- <= FPGA_IN_pHOLD-;
END IF;
END PROCESS;



VGA_RAM_READ_DATA <= NOT(SYNTHESIZED_WIRE_262 OR SYNTHESIZED_WIRE_263);


PROCESS(SYNTHESIZED_WIRE_265,SYNTHESIZED_WIRE_264,SYNTHESIZED_WIRE_674)
BEGIN
IF (SYNTHESIZED_WIRE_264 = '0') THEN
	PS2_KEYBOARD_STATUS <= '0';
ELSIF (SYNTHESIZED_WIRE_674 = '0') THEN
	PS2_KEYBOARD_STATUS <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_265)) THEN
	PS2_KEYBOARD_STATUS <= SYNTHESIZED_WIRE_674;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_309 <= NOT(OUT_sMEMR);



SYNTHESIZED_WIRE_94 <= NOT(READ_RAM);



SYNTHESIZED_WIRE_722 <= FPGA_ROM- AND SYNTHESIZED_WIRE_665 AND Z80_MREQ AND Z80_MREQ;


SYNTHESIZED_WIRE_0 <= FPGA_IN_XRDY AND FPGA_IN_RDY AND BOARD_WAIT-;


Z80_WR <= NOT(Z80_WR-);



SYNTHESIZED_WIRE_721 <= NOT(PORT_SELECT_6C- OR OUT_pWR-);


ROM_OE <= SYNTHESIZED_WIRE_269 AND OUT_pDBIN AND FPGA_ROM;


SYNTHESIZED_WIRE_262 <= NOT(OUT_sMEMR AND VGA_RAM_SELECT);


SYNTHESIZED_WIRE_263 <= NOT(OUT_pDBIN);




ROM_ADDRESS(5) <= S100_A5 OR S100_A5;


ROM_ADDRESS(4) <= S100_A4 OR S100_A4;


ROM_ADDRESS(3) <= S100_A3 OR S100_A3;


ROM_ADDRESS(2) <= S100_A2 OR S100_A2;


ROM_ADDRESS(1) <= S100_A1 OR S100_A1;


Z80_IORQ <= NOT(Z80_IORQ-);



ROM_ADDRESS(0) <= S100_A0 OR S100_A0;


ROM_ADDRESS(11) <= S100_A11 OR S100_A11;


ROM_ADDRESS(10) <= S100_A10 OR S100_A10;


ROM_ADDRESS(9) <= S100_A9 OR S100_A9;


ROM_ADDRESS(8) <= S100_A8 OR S100_A8;


ROM_ADDRESS(7) <= S100_A7 OR S100_A7;


ROM_ADDRESS(6) <= S100_A6 OR S100_A6;


ROM_ADDRESS(12) <= ROM_A12 OR ROM_A12;


FPGA_ROM <= NOT(FPGA_ROM-);



VGA_RAM_SELECT <= NOT(SYNTHESIZED_WIRE_270);



Z80_RD <= NOT(Z80_RD-);




b2v_inst321 : 74684_20
PORT MAP(P2 => SYNTHESIZED_WIRE_675,
		 Q2 => SYNTHESIZED_WIRE_675,
		 P1 => SYNTHESIZED_WIRE_675,
		 Q1 => SYNTHESIZED_WIRE_675,
		 P0 => SYNTHESIZED_WIRE_675,
		 Q0 => SYNTHESIZED_WIRE_675,
		 P7 => S100_A15,
		 Q7 => SYNTHESIZED_WIRE_676,
		 Q6 => SYNTHESIZED_WIRE_676,
		 P6 => S100_A14,
		 Q5 => SYNTHESIZED_WIRE_676,
		 P5 => S100_A13,
		 P4 => S100_A12,
		 Q4 => SYNTHESIZED_WIRE_675,
		 Q3 => SYNTHESIZED_WIRE_675,
		 P3 => SYNTHESIZED_WIRE_675,
		 EQUALN => SYNTHESIZED_WIRE_270);


S100_PHANTOM_LED <= NOT(SYNTHESIZED_WIRE_283);



VGA_RAM_READ_DATA- <= NOT(VGA_RAM_READ_DATA);




PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_285,SYNTHESIZED_WIRE_284,Z80_LOCAL_D0)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	CTL <= '0';
ELSIF (SYNTHESIZED_WIRE_285 = '0') THEN
	CTL <= '1';
ELSIF (SYNTHESIZED_WIRE_284 = '1') THEN
	CTL <= Z80_LOCAL_D0;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_286 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_269 <= NOT(pSYNC_RAW);



SYNTHESIZED_WIRE_284 <= NOT(OUT_pWR- OR SYNTHESIZED_WIRE_286 OR PORT_C2H-);


SYNTHESIZED_WIRE_67 <= NOT(SYNTHESIZED_WIRE_677);



Z80_MREQ <= NOT(Z80_MREQ-);



SYNTHESIZED_WIRE_660 <= NOT(OUT_pDBIN);



b2v_inst331 : 74373b_21
PORT MAP(G => SYNTHESIZED_WIRE_660,
		 OEN => SYNTHESIZED_WIRE_678,
		 D => CURSOR_Y,
		 Q => Z80_LOCAL_DI);


VGA_CURSOR_OE- <= SYNTHESIZED_WIRE_668 AND SYNTHESIZED_WIRE_669 AND SYNTHESIZED_WIRE_678;


b2v_inst333 : 74138_22
PORT MAP(A => S100_A0,
		 B => S100_A1,
		 G1 => SYNTHESIZED_WIRE_293,
		 C => SYNTHESIZED_WIRE_294,
		 G2AN => SYNTHESIZED_WIRE_679,
		 G2BN => SYNTHESIZED_WIRE_679,
		 Y0N => PORT_SELECT_68-,
		 Y1N => PORT_SELECT_69-,
		 Y2N => PORT_SELECT_6A-,
		 Y3N => PORT_SELECT_6B-);


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_659,SYNTHESIZED_WIRE_297,Z80_LOCAL_D0(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	FPGA_OUT_PRN_STROBE <= '0';
ELSIF (SYNTHESIZED_WIRE_659 = '0') THEN
	FPGA_OUT_PRN_STROBE <= '1';
ELSIF (SYNTHESIZED_WIRE_297 = '1') THEN
	FPGA_OUT_PRN_STROBE <= Z80_LOCAL_D0;
END IF;
END PROCESS;


b2v_inst335 : 74244_23
PORT MAP(1A2 => FPGA_IN_PRN_BUSY,
		 1A4 => SYNTHESIZED_WIRE_680,
		 1A1 => DFF_inst143,
		 1A3 => SYNTHESIZED_WIRE_680,
		 1GN => PRINTER_STATUS_PORT-,
		 2A3 => SYNTHESIZED_WIRE_680,
		 2GN => PRINTER_STATUS_PORT-,
		 2A1 => SYNTHESIZED_WIRE_680,
		 2A4 => SYNTHESIZED_WIRE_680,
		 2A2 => SYNTHESIZED_WIRE_680,
		 1Y2 => Z80_LOCAL_DI(1),
		 1Y4 => Z80_LOCAL_DI(3),
		 2Y1 => Z80_LOCAL_DI(4),
		 1Y1 => Z80_LOCAL_DI(0),
		 2Y3 => Z80_LOCAL_DI(6),
		 2Y4 => Z80_LOCAL_DI(7),
		 1Y3 => Z80_LOCAL_DI(2),
		 2Y2 => Z80_LOCAL_DI(5));


PROCESS(SYNTHESIZED_WIRE_305,IN_BOARD_RESET-,SYNTHESIZED_WIRE_306)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DFF_inst336 <= '0';
ELSIF (SYNTHESIZED_WIRE_306 = '0') THEN
	DFF_inst336 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_305)) THEN
	DFF_inst336 <= Z80_LOCAL_D0(7);
END IF;
END PROCESS;



SYNTHESIZED_WIRE_95 <= NOT(OUT_sOUT);



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_671,PS2_DATA_IN,SYNTHESIZED_WIRE_307)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_154 <= '0';
ELSIF (SYNTHESIZED_WIRE_671 = '0') THEN
	SYNTHESIZED_WIRE_154 <= '1';
ELSIF (PS2_DATA_IN = '1') THEN
	SYNTHESIZED_WIRE_154 <= SYNTHESIZED_WIRE_307;
END IF;
END PROCESS;


FPGA_ROM- <= SYNTHESIZED_WIRE_309 OR DISABLE_ALL_ROM OR SYNTHESIZED_WIRE_665;


SYNTHESIZED_WIRE_311 <= NOT(OUT_pDBIN);



PS2_DATA_IN <= NOT(PS2_DATA- OR SYNTHESIZED_WIRE_311);


FORCE_LOW_SPEED- <= NOT(DFF_inst336);



SYNTHESIZED_WIRE_316 <= SPI_READ OR SPI_WRITE;


BUZZER <= NOT(START_BUZZER);



PROCESS(SYNTHESIZED_WIRE_313,SYNTHESIZED_WIRE_681,SYNTHESIZED_WIRE_682)
BEGIN
IF (SYNTHESIZED_WIRE_681 = '0') THEN
	START_BUZZER <= '0';
ELSIF (SYNTHESIZED_WIRE_682 = '0') THEN
	START_BUZZER <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_313)) THEN
	START_BUZZER <= SYNTHESIZED_WIRE_682;
END IF;
END PROCESS;


F_BOARD_ACTIVE- <= SYNTHESIZED_WIRE_683 AND CPU_CLK_COUNTER(20);


b2v_inst347 : spi_16bit_master
GENERIC MAP(d_width => 16,
			slaves => 4
			)
PORT MAP(clock => SPI_CLK,
		 reset_n => IN_BOARD_RESET-,
		 enable => SYNTHESIZED_WIRE_316,
		 cpol => SYNTHESIZED_WIRE_684,
		 cpha => SYNTHESIZED_WIRE_684,
		 cont => SYNTHESIZED_WIRE_319,
		 miso => RTC_SPI_SO,
		 addr => SPI_INPUT_CS,
		 clk_div => SPI_CLK_DIV,
		 tx_data => SPI_DATA_OUT_BUS,
		 sclk => SPI_MASTER_CLK,
		 mosi => RTC_SPI_SI,
		 busy => SPI_BUSY_FLAG,
		 rx_data => SPI_DATA_IN_BUS);


SYNTHESIZED_WIRE_658 <= NOT(OUT_pWR- OR SYNTHESIZED_WIRE_320 OR PORT_C7H-);


PROCESS(COUNTER_BUS(16),SYNTHESIZED_WIRE_681,SYNTHESIZED_WIRE_322)
BEGIN
IF (SYNTHESIZED_WIRE_681 = '0') THEN
	DFF_inst349 <= '0';
ELSIF (SYNTHESIZED_WIRE_322 = '0') THEN
	DFF_inst349 <= '1';
ELSIF (RISING_EDGE(COUNTER_BUS(16))) THEN
	DFF_inst349 <= START_BUZZER;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_589 <= NOT(Z80_HALT-);




PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_323,PS2_STATUS_IN,PS2_KEYBOARD_STATUS)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_107 <= '0';
ELSIF (SYNTHESIZED_WIRE_323 = '0') THEN
	SYNTHESIZED_WIRE_107 <= '1';
ELSIF (PS2_STATUS_IN = '1') THEN
	SYNTHESIZED_WIRE_107 <= PS2_KEYBOARD_STATUS;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_324 <= NOT(OUT_pDBIN);



PS2_STATUS_IN <= NOT(PS2_STATUS- OR SYNTHESIZED_WIRE_324);




SYNTHESIZED_WIRE_320 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_297 <= NOT(OUT_pWR- OR SYNTHESIZED_WIRE_325 OR PORT_C6H-);


PROCESS(COUNTER_BUS(16),SYNTHESIZED_WIRE_681,SYNTHESIZED_WIRE_327)
BEGIN
IF (SYNTHESIZED_WIRE_681 = '0') THEN
	DFF_inst358 <= '0';
ELSIF (SYNTHESIZED_WIRE_327 = '0') THEN
	DFF_inst358 <= '1';
ELSIF (RISING_EDGE(COUNTER_BUS(16))) THEN
	DFF_inst358 <= DFF_inst349;
END IF;
END PROCESS;


PRINTER_STATUS_PORT- <= NOT(OUT_pDBIN AND OUT_sINP AND SYNTHESIZED_WIRE_328);


Z80_M1 <= NOT(Z80_M1-);



SYNTHESIZED_WIRE_328 <= NOT(PORT_C7H-);




STOP_BUZZER <= NOT(DFF_inst358);



SYNTHESIZED_WIRE_325 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_681 <= IN_BOARD_RESET- AND STOP_BUZZER;


SYNTHESIZED_WIRE_70 <= NOT(SYNTHESIZED_WIRE_658);




SYNTHESIZED_WIRE_313 <= NOT(OUT_pWR- OR SYNTHESIZED_WIRE_330 OR PORT_0-);


SYNTHESIZED_WIRE_330 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_351 <= NOT(PORT_SELECT_6B- OR OUT_pWR-);


b2v_inst37 : 74164_24
PORT MAP(CLRN => SYNTHESIZED_WIRE_331,
		 CLK => OUT_CPU_CLK,
		 B => SYNTHESIZED_WIRE_332,
		 A => USB_DATA_OUT,
		 QB => SYNTHESIZED_WIRE_606);


SYNTHESIZED_WIRE_372 <= NOT(PORT_SELECT_6B- OR SYNTHESIZED_WIRE_333);



SPI_CLK_DIV <= NOT(SYNTHESIZED_WIRE_685);




SPI_INPUT_CS <= NOT(SYNTHESIZED_WIRE_685);



b2v_inst375 : 74148_25
PORT MAP(5N => SYNTHESIZED_WIRE_336,
		 0N => SYNTHESIZED_WIRE_337,
		 1N => SYNTHESIZED_WIRE_338,
		 2N => SYNTHESIZED_WIRE_339,
		 3N => SYNTHESIZED_WIRE_340,
		 4N => SYNTHESIZED_WIRE_341,
		 EIN => SYNTHESIZED_WIRE_342,
		 6N => SYNTHESIZED_WIRE_343,
		 7N => SYNTHESIZED_WIRE_344,
		 A1N => SYNTHESIZED_WIRE_481,
		 A0N => SYNTHESIZED_WIRE_479,
		 A2N => SYNTHESIZED_WIRE_484,
		 GSN => SYNTHESIZED_WIRE_482);


b2v_inst376 : 74373_26
PORT MAP(D1 => SYNTHESIZED_WIRE_686,
		 D3 => RTC_INT,
		 D6 => FPGA_IN_INT_B-,
		 D7 => FPGA_IN_INT_A-,
		 D2 => SYNTHESIZED_WIRE_686,
		 G => SYNTHESIZED_WIRE_687,
		 D4 => FPGA_IN_INT_D-,
		 D5 => FPGA_IN_INT_C-,
		 D8 => SYNTHESIZED_WIRE_686,
		 OEN => SYNTHESIZED_WIRE_349,
		 Q3 => SYNTHESIZED_WIRE_340,
		 Q6 => SYNTHESIZED_WIRE_343,
		 Q7 => SYNTHESIZED_WIRE_344,
		 Q2 => SYNTHESIZED_WIRE_339,
		 Q8 => SYNTHESIZED_WIRE_337,
		 Q4 => SYNTHESIZED_WIRE_341,
		 Q5 => SYNTHESIZED_WIRE_336,
		 Q1 => SYNTHESIZED_WIRE_338);


PROCESS(SYNTHESIZED_WIRE_351,SYNTHESIZED_WIRE_688,SYNTHESIZED_WIRE_689)
BEGIN
IF (SYNTHESIZED_WIRE_688 = '0') THEN
	DFF_inst377 <= '0';
ELSIF (SYNTHESIZED_WIRE_689 = '0') THEN
	DFF_inst377 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_351)) THEN
	DFF_inst377 <= SYNTHESIZED_WIRE_689;
END IF;
END PROCESS;



PROCESS(SPI_CLK,SYNTHESIZED_WIRE_688,SYNTHESIZED_WIRE_689)
BEGIN
IF (SYNTHESIZED_WIRE_688 = '0') THEN
	SPI_WRITE <= '0';
ELSIF (SYNTHESIZED_WIRE_689 = '0') THEN
	SPI_WRITE <= '1';
ELSIF (RISING_EDGE(SPI_CLK)) THEN
	SPI_WRITE <= DFF_inst377;
END IF;
END PROCESS;


DATA_OUT_D6 <= Z80_LOCAL_D0(6) OR Z80_LOCAL_D0(6);


SYNTHESIZED_WIRE_356 <= NOT(SPI_BUSY_FLAG);



SYNTHESIZED_WIRE_688 <= SYNTHESIZED_WIRE_356 AND IN_BOARD_RESET-;


SPI_CLK <= NOT(COUNTER_BUS(4));




SYNTHESIZED_WIRE_333 <= NOT(OUT_pDBIN);



b2v_inst385 : 74138_27
PORT MAP(A => S100_A0,
		 B => S100_A1,
		 G1 => SYNTHESIZED_WIRE_357,
		 C => SYNTHESIZED_WIRE_358,
		 G2AN => SYNTHESIZED_WIRE_690,
		 G2BN => SYNTHESIZED_WIRE_690,
		 Y0N => PORT_SELECT_6C-,
		 Y1N => PORT_SELECT_6D-,
		 Y2N => PORT_SELECT_6E-,
		 Y3N => PORT_SELECT_6F-);


b2v_inst386 : 74684_28
PORT MAP(P2 => S100_A2,
		 Q2 => SYNTHESIZED_WIRE_691,
		 P1 => SYNTHESIZED_WIRE_691,
		 Q1 => SYNTHESIZED_WIRE_691,
		 P0 => SYNTHESIZED_WIRE_691,
		 Q0 => SYNTHESIZED_WIRE_691,
		 P7 => S100_A7,
		 Q7 => SYNTHESIZED_WIRE_691,
		 Q6 => SYNTHESIZED_WIRE_692,
		 P6 => S100_A6,
		 Q5 => SYNTHESIZED_WIRE_692,
		 P5 => S100_A5,
		 P4 => S100_A4,
		 Q4 => SYNTHESIZED_WIRE_691,
		 Q3 => SYNTHESIZED_WIRE_692,
		 P3 => S100_A3,
		 EQUALN => SYNTHESIZED_WIRE_679);


PROCESS(SYNTHESIZED_WIRE_372,SYNTHESIZED_WIRE_693,SYNTHESIZED_WIRE_694)
BEGIN
IF (SYNTHESIZED_WIRE_693 = '0') THEN
	DFF_inst387 <= '0';
ELSIF (SYNTHESIZED_WIRE_694 = '0') THEN
	DFF_inst387 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_372)) THEN
	DFF_inst387 <= SYNTHESIZED_WIRE_694;
END IF;
END PROCESS;



PROCESS(SPI_CLK,SYNTHESIZED_WIRE_693,SYNTHESIZED_WIRE_694)
BEGIN
IF (SYNTHESIZED_WIRE_693 = '0') THEN
	SPI_READ <= '0';
ELSIF (SYNTHESIZED_WIRE_694 = '0') THEN
	SPI_READ <= '1';
ELSIF (RISING_EDGE(SPI_CLK)) THEN
	SPI_READ <= DFF_inst387;
END IF;
END PROCESS;


DATA_OUT_D7 <= Z80_LOCAL_D0(7) OR Z80_LOCAL_D0(7);


SYNTHESIZED_WIRE_377 <= NOT(SPI_BUSY_FLAG);



SYNTHESIZED_WIRE_693 <= SYNTHESIZED_WIRE_377 AND IN_BOARD_RESET-;


SYNTHESIZED_WIRE_704 <= NOT(OUT_pWR- OR PORT_SELECT_68- OR SYNTHESIZED_WIRE_378);




SYNTHESIZED_WIRE_293 <= OUT_sINP OR OUT_sOUT;


SYNTHESIZED_WIRE_378 <= NOT(OUT_sOUT);



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_379,Z80_LOCAL_D0(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	RTC_CS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	RTC_CS <= '1';
ELSIF (SYNTHESIZED_WIRE_379 = '1') THEN
	RTC_CS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_379 <= NOT(OUT_pWR- OR PORT_SELECT_6A- OR SYNTHESIZED_WIRE_381);


SYNTHESIZED_WIRE_381 <= NOT(OUT_sOUT);



b2v_inst4 : pll01_50
PORT MAP(inclk0 => 50mHz,
		 c0 => 2mHz,
		 c1 => 400_KHz_CLK,
		 c2 => 10mHz,
		 c3 => 25Mhz);





PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(7))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_7_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_7_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_7_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(6))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_6_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_6_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_6_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(5))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_5_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_5_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_5_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(4))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_4_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_4_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_4_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(3))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_3_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_3_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_3_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(2))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_2_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_2_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_2_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(1))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_1_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_1_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_1_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_696,SPI_DATA_IN_BUS(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_IN_0_A <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	DATA_IN_0_A <= '1';
ELSIF (SYNTHESIZED_WIRE_696 = '1') THEN
	DATA_IN_0_A <= SPI_DATA_IN_BUS;
END IF;
END PROCESS;


READ_RAM <= NOT(OUT_RAM_READ-);



b2v_inst410 : 74244_29
PORT MAP(1A2 => DATA_IN_6_A,
		 1A4 => DATA_IN_4_A,
		 1A1 => DATA_IN_7_A,
		 1A3 => DATA_IN_5_A,
		 1GN => SYNTHESIZED_WIRE_698,
		 2A3 => DATA_IN_1_A,
		 2GN => SYNTHESIZED_WIRE_698,
		 2A1 => DATA_IN_3_A,
		 2A4 => DATA_IN_0_A,
		 2A2 => DATA_IN_2_A,
		 1Y2 => Z80_LOCAL_DI(6),
		 1Y4 => Z80_LOCAL_DI(4),
		 2Y1 => Z80_LOCAL_DI(3),
		 1Y1 => Z80_LOCAL_DI(7),
		 2Y3 => Z80_LOCAL_DI(1),
		 2Y4 => Z80_LOCAL_DI(0),
		 1Y3 => Z80_LOCAL_DI(5),
		 2Y2 => Z80_LOCAL_DI(2));


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_697,SYNTHESIZED_WIRE_699,SPI_BUSY_FLAG)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_702 <= '0';
ELSIF (SYNTHESIZED_WIRE_697 = '0') THEN
	SYNTHESIZED_WIRE_702 <= '1';
ELSIF (SYNTHESIZED_WIRE_699 = '1') THEN
	SYNTHESIZED_WIRE_702 <= SPI_BUSY_FLAG;
END IF;
END PROCESS;


b2v_inst412 : 74684_30
PORT MAP(P2 => S100_A2,
		 Q2 => SYNTHESIZED_WIRE_700,
		 P1 => SYNTHESIZED_WIRE_701,
		 Q1 => SYNTHESIZED_WIRE_701,
		 P0 => SYNTHESIZED_WIRE_701,
		 Q0 => SYNTHESIZED_WIRE_701,
		 P7 => S100_A7,
		 Q7 => SYNTHESIZED_WIRE_701,
		 Q6 => SYNTHESIZED_WIRE_700,
		 P6 => S100_A6,
		 Q5 => SYNTHESIZED_WIRE_700,
		 P5 => S100_A5,
		 P4 => S100_A4,
		 Q4 => SYNTHESIZED_WIRE_701,
		 Q3 => SYNTHESIZED_WIRE_700,
		 P3 => S100_A3,
		 EQUALN => SYNTHESIZED_WIRE_690);


b2v_inst413 : 74244_31
PORT MAP(1A2 => SYNTHESIZED_WIRE_702,
		 1A4 => SYNTHESIZED_WIRE_702,
		 1A1 => SYNTHESIZED_WIRE_702,
		 1A3 => SYNTHESIZED_WIRE_702,
		 1GN => SYNTHESIZED_WIRE_703,
		 2A3 => SYNTHESIZED_WIRE_702,
		 2GN => SYNTHESIZED_WIRE_703,
		 2A1 => SYNTHESIZED_WIRE_702,
		 2A4 => SYNTHESIZED_WIRE_702,
		 2A2 => SYNTHESIZED_WIRE_702,
		 1Y2 => Z80_LOCAL_DI(6),
		 1Y4 => Z80_LOCAL_DI(4),
		 2Y1 => Z80_LOCAL_DI(3),
		 1Y1 => Z80_LOCAL_DI(7),
		 2Y3 => Z80_LOCAL_DI(1),
		 2Y4 => Z80_LOCAL_DI(0),
		 1Y3 => Z80_LOCAL_DI(5),
		 2Y2 => Z80_LOCAL_DI(2));


SYNTHESIZED_WIRE_696 <= OUT_pDBIN AND SYNTHESIZED_WIRE_422 AND OUT_sINP;


SYNTHESIZED_WIRE_422 <= NOT(PORT_SELECT_69-);



SPI_RTC_READ_DATA- <= NOT(SYNTHESIZED_WIRE_696 OR SYNTHESIZED_WIRE_699);


SYNTHESIZED_WIRE_698 <= NOT(SYNTHESIZED_WIRE_696);



SYNTHESIZED_WIRE_699 <= OUT_pDBIN AND SYNTHESIZED_WIRE_426 AND OUT_sINP;


SYNTHESIZED_WIRE_426 <= NOT(PORT_SELECT_6A-);



SYNTHESIZED_WIRE_245 <= NOT(SYNTHESIZED_WIRE_427 OR OUT_pWR- OR PORT_7-);


SYNTHESIZED_WIRE_703 <= NOT(SYNTHESIZED_WIRE_699);




PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(7))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(6))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(5))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(4))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(3))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(2))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(1))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_695,SYNTHESIZED_WIRE_704,Z80_LOCAL_D0(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_695 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_704 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_243 <= NOT(SYNTHESIZED_WIRE_445 OR OUT_pWR- OR PORT_7-);


SYNTHESIZED_WIRE_92 <= VGA_RAM_READ_DATA- AND VGA_CURSOR_OE- AND SPI_RTC_READ_DATA-;



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(7))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(6))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(5))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(4))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(3))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(2))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(1))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_706,SYNTHESIZED_WIRE_705,Z80_LOCAL_D0(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_DATA_OUT_BUS <= '0';
ELSIF (SYNTHESIZED_WIRE_706 = '0') THEN
	SPI_DATA_OUT_BUS <= '1';
ELSIF (SYNTHESIZED_WIRE_705 = '1') THEN
	SPI_DATA_OUT_BUS <= Z80_LOCAL_D0;
END IF;
END PROCESS;


b2v_inst44 : fpga_rom_16k
PORT MAP(clock => ROM_OE,
		 address => ROM_ADDRESS,
		 q => SYNTHESIZED_WIRE_604);


SYNTHESIZED_WIRE_705 <= NOT(OUT_pWR- OR PORT_SELECT_69- OR SYNTHESIZED_WIRE_462);


SYNTHESIZED_WIRE_462 <= NOT(OUT_sOUT);





SYNTHESIZED_WIRE_464 <= NOT(SYNTHESIZED_WIRE_687);



SYNTHESIZED_WIRE_465 <= NOT(SYNTHESIZED_WIRE_464);



SYNTHESIZED_WIRE_466 <= NOT(SYNTHESIZED_WIRE_465);



SYNTHESIZED_WIRE_467 <= NOT(SYNTHESIZED_WIRE_466);



SYNTHESIZED_WIRE_468 <= NOT(SYNTHESIZED_WIRE_467);



SYNTHESIZED_WIRE_469 <= NOT(SYNTHESIZED_WIRE_468);



PROCESS(DATA_OUT_D0,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D0 <= DATA_OUT_D0;
ELSE
	FPGA_BI_D0 <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_470 <= NOT(SYNTHESIZED_WIRE_469);



SYNTHESIZED_WIRE_483 <= NOT(SYNTHESIZED_WIRE_470);



b2v_inst452 : 74244_32
PORT MAP(1A2 => SYNTHESIZED_WIRE_707,
		 1A4 => SYNTHESIZED_WIRE_472,
		 1A1 => SYNTHESIZED_WIRE_707,
		 1A3 => SYNTHESIZED_WIRE_707,
		 1GN => INTA_READ_DATA-,
		 2A3 => SYNTHESIZED_WIRE_707,
		 2GN => INTA_READ_DATA-,
		 2A1 => SYNTHESIZED_WIRE_476,
		 2A4 => SYNTHESIZED_WIRE_707,
		 2A2 => SYNTHESIZED_WIRE_478,
		 1Y2 => Z80_LOCAL_DI(1),
		 1Y4 => Z80_LOCAL_DI(3),
		 2Y1 => Z80_LOCAL_DI(4),
		 1Y1 => Z80_LOCAL_DI(0),
		 2Y3 => Z80_LOCAL_DI(6),
		 2Y4 => Z80_LOCAL_DI(7),
		 1Y3 => Z80_LOCAL_DI(2),
		 2Y2 => Z80_LOCAL_DI(5));


SYNTHESIZED_WIRE_472 <= NOT(SYNTHESIZED_WIRE_479);



SYNTHESIZED_WIRE_93 <= PRINTER_STATUS_PORT- AND INTA_READ_DATA-;


BOARD_INT- <= SYNTHESIZED_WIRE_480 AND S100_INT-;


SYNTHESIZED_WIRE_687 <= NOT(OUT_sINTA);



SYNTHESIZED_WIRE_476 <= NOT(SYNTHESIZED_WIRE_481);



SYNTHESIZED_WIRE_480 <= FPGA_IN_ENABLE_INTA OR SYNTHESIZED_WIRE_482;


INTA_READ_DATA- <= SYNTHESIZED_WIRE_483 OR FPGA_IN_ENABLE_INTA;


PROCESS(FPGA_BI_D0,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(0) <= FPGA_BI_D0;
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;




SYNTHESIZED_WIRE_478 <= NOT(SYNTHESIZED_WIRE_484);




SYNTHESIZED_WIRE_357 <= OUT_sINP OR OUT_sOUT;


SYNTHESIZED_WIRE_511 <= NOT(PORT_SELECT_6D- OR OUT_pWR-);



SYNTHESIZED_WIRE_723 <= NOT(PORT_SELECT_6E- OR OUT_pWR-);


PROCESS(SYNTHESIZED_WIRE_486,SYNTHESIZED_WIRE_708,SYNTHESIZED_WIRE_709)
BEGIN
IF (SYNTHESIZED_WIRE_708 = '0') THEN
	DFF_inst468 <= '0';
ELSIF (SYNTHESIZED_WIRE_709 = '0') THEN
	DFF_inst468 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_486)) THEN
	DFF_inst468 <= SYNTHESIZED_WIRE_709;
END IF;
END PROCESS;


b2v_inst469 : 74244_33
PORT MAP(1A2 => SDCARD_OUT_6,
		 1A4 => SDCARD_OUT_4,
		 1A1 => SDCARD_OUT_7,
		 1A3 => SDCARD_OUT_5,
		 1GN => SYNTHESIZED_WIRE_710,
		 2A3 => SDCARD_OUT_1,
		 2GN => SYNTHESIZED_WIRE_710,
		 2A1 => SDCARD_OUT_3,
		 2A4 => SDCARD_OUT_0,
		 2A2 => SDCARD_OUT_2,
		 1Y2 => Z80_LOCAL_DI(6),
		 1Y4 => Z80_LOCAL_DI(4),
		 2Y1 => Z80_LOCAL_DI(3),
		 1Y1 => Z80_LOCAL_DI(7),
		 2Y3 => Z80_LOCAL_DI(1),
		 2Y4 => Z80_LOCAL_DI(0),
		 1Y3 => Z80_LOCAL_DI(5),
		 2Y2 => Z80_LOCAL_DI(2));


PROCESS(DATA_OUT_D1,WRITE_RAM)
BEGIN
if (WRITE_RAM = '1') THEN
	FPGA_BI_D1 <= DATA_OUT_D1;
ELSE
	FPGA_BI_D1 <= 'Z';
END IF;
END PROCESS;


SD_CARD_READ_DATA- <= NOT(SYNTHESIZED_WIRE_711 OR SYNTHESIZED_WIRE_712);


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_712,SD_CARD_BUSY)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_497 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SYNTHESIZED_WIRE_497 <= '1';
ELSIF (SYNTHESIZED_WIRE_712 = '1') THEN
	SYNTHESIZED_WIRE_497 <= SD_CARD_BUSY;
END IF;
END PROCESS;


b2v_inst472 : 74244_34
PORT MAP(1A2 => SYNTHESIZED_WIRE_714,
		 1A4 => SYNTHESIZED_WIRE_714,
		 1A1 => SYNTHESIZED_WIRE_497,
		 1A3 => SYNTHESIZED_WIRE_714,
		 1GN => SYNTHESIZED_WIRE_715,
		 2A3 => SYNTHESIZED_WIRE_500,
		 2GN => SYNTHESIZED_WIRE_715,
		 2A1 => SYNTHESIZED_WIRE_714,
		 2A4 => SYNTHESIZED_WIRE_503,
		 2A2 => SYNTHESIZED_WIRE_714,
		 1Y2 => Z80_LOCAL_DI(6),
		 1Y4 => Z80_LOCAL_DI(4),
		 2Y1 => Z80_LOCAL_DI(3),
		 1Y1 => Z80_LOCAL_DI(7),
		 2Y3 => Z80_LOCAL_DI(1),
		 2Y4 => Z80_LOCAL_DI(0),
		 1Y3 => Z80_LOCAL_DI(5),
		 2Y2 => Z80_LOCAL_DI(2));


SYNTHESIZED_WIRE_711 <= OUT_pDBIN AND SYNTHESIZED_WIRE_505;


SYNTHESIZED_WIRE_712 <= OUT_pDBIN AND SYNTHESIZED_WIRE_506;


SYNTHESIZED_WIRE_715 <= NOT(SYNTHESIZED_WIRE_712);



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_712,SYNTHESIZED_WIRE_716)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_500 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SYNTHESIZED_WIRE_500 <= '1';
ELSIF (SYNTHESIZED_WIRE_712 = '1') THEN
	SYNTHESIZED_WIRE_500 <= SYNTHESIZED_WIRE_716;
END IF;
END PROCESS;



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_511,Z80_LOCAL_D0(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SPI_SD_CLK_SPEED <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	SPI_SD_CLK_SPEED <= '1';
ELSIF (SYNTHESIZED_WIRE_511 = '1') THEN
	SPI_SD_CLK_SPEED <= Z80_LOCAL_D0;
END IF;
END PROCESS;


b2v_inst479 : 21mux_35
PORT MAP(S => SPI_SD_CLK_SPEED,
		 B => 400_KHz_CLK,
		 A => 10mHz,
		 Y => LOCAL_SD_SPI_CLK);


b2v_inst48 : 74138_36
PORT MAP(A => S100_A0,
		 B => S100_A1,
		 G1 => SYNTHESIZED_WIRE_513,
		 C => S100_A2,
		 G2AN => SYNTHESIZED_WIRE_718,
		 G2BN => SYNTHESIZED_WIRE_718,
		 Y0N => PORT_C0H-,
		 Y1N => PORT_C1H-,
		 Y2N => PORT_C2H-,
		 Y6N => PORT_C6H-,
		 Y7N => PORT_C7H-);


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_712,SYNTHESIZED_WIRE_719)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_503 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SYNTHESIZED_WIRE_503 <= '1';
ELSIF (SYNTHESIZED_WIRE_712 = '1') THEN
	SYNTHESIZED_WIRE_503 <= SYNTHESIZED_WIRE_719;
END IF;
END PROCESS;



PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(7))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_7 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_7 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_7 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(6))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_6 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_6 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_6 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(5))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_5 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_5 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_5 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(4))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_4 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_4 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_4 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(3))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_3 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_3 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_3 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(2))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_2 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_2 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_2 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(1))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_1 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_1 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_1 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_713,SYNTHESIZED_WIRE_711,DATA_FROM_SDCARD(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	SDCARD_OUT_0 <= '0';
ELSIF (SYNTHESIZED_WIRE_713 = '0') THEN
	SDCARD_OUT_0 <= '1';
ELSIF (SYNTHESIZED_WIRE_711 = '1') THEN
	SDCARD_OUT_0 <= DATA_FROM_SDCARD;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_605 <= NOT(IN_BOARD_RESET-);



b2v_inst490 : spi_master
GENERIC MAP(d_width => 8,
			slaves => 2
			)
PORT MAP(clock => LOCAL_SD_SPI_CLK,
		 reset_n => IN_BOARD_RESET-,
		 enable => SYNTHESIZED_WIRE_535,
		 cpol => SYNTHESIZED_WIRE_720,
		 cpha => SYNTHESIZED_WIRE_720,
		 cont => SYNTHESIZED_WIRE_720,
		 miso => SD_DO,
		 addr => SD_CARD_ADDRESS,
		 clk_div => SD_CARD_CLK_DIV,
		 tx_data => DATA_TO_SDCARD,
		 sclk => SD_CLK,
		 mosi => SD_CMD,
		 busy => SD_CARD_BUSY,
		 rx_data => DATA_FROM_SDCARD,
		 ss_n => SD_SLAVES);


SYNTHESIZED_WIRE_505 <= NOT(PORT_SELECT_6C-);



SYNTHESIZED_WIRE_506 <= NOT(PORT_SELECT_6E-);



SYNTHESIZED_WIRE_710 <= NOT(SYNTHESIZED_WIRE_711);




PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(7))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(6))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(5))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(4))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(3))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;


b2v_inst5 : counter01_32
PORT MAP(clock => 2mHz,
		 q => COUNTER_BUS);


OUT_RAM_READ- <= NOT(MEM_READ AND SYNTHESIZED_WIRE_722);


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(2))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(1))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(IN_BOARD_RESET-,SYNTHESIZED_WIRE_717,SYNTHESIZED_WIRE_721,Z80_LOCAL_D0(0))
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	DATA_TO_SDCARD <= '0';
ELSIF (SYNTHESIZED_WIRE_717 = '0') THEN
	DATA_TO_SDCARD <= '1';
ELSIF (SYNTHESIZED_WIRE_721 = '1') THEN
	DATA_TO_SDCARD <= Z80_LOCAL_D0;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_535 <= SD_READ OR SD_WRITE;



PROCESS(LOCAL_SD_SPI_CLK,SYNTHESIZED_WIRE_708,SYNTHESIZED_WIRE_709)
BEGIN
IF (SYNTHESIZED_WIRE_708 = '0') THEN
	SD_WRITE <= '0';
ELSIF (SYNTHESIZED_WIRE_709 = '0') THEN
	SD_WRITE <= '1';
ELSIF (RISING_EDGE(LOCAL_SD_SPI_CLK)) THEN
	SD_WRITE <= DFF_inst468;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_708 <= SYNTHESIZED_WIRE_559 AND IN_BOARD_RESET-;


PROCESS(SYNTHESIZED_WIRE_717,IN_BOARD_RESET-,SYNTHESIZED_WIRE_723,Z80_LOCAL_D0(0))
BEGIN
IF (SYNTHESIZED_WIRE_717 = '0') THEN
	SYNTHESIZED_WIRE_716 <= '0';
ELSIF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_716 <= '1';
ELSIF (SYNTHESIZED_WIRE_723 = '1') THEN
	SYNTHESIZED_WIRE_716 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_717,IN_BOARD_RESET-,SYNTHESIZED_WIRE_723,Z80_LOCAL_D0(1))
BEGIN
IF (SYNTHESIZED_WIRE_717 = '0') THEN
	SYNTHESIZED_WIRE_719 <= '0';
ELSIF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_719 <= '1';
ELSIF (SYNTHESIZED_WIRE_723 = '1') THEN
	SYNTHESIZED_WIRE_719 <= Z80_LOCAL_D0;
END IF;
END PROCESS;


PROCESS(FPGA_BI_D1,READ_RAM)
BEGIN
if (READ_RAM = '1') THEN
	Z80_LOCAL_DI(1) <= FPGA_BI_D1;
ELSE
	Z80_LOCAL_DI(1) <= 'Z';
END IF;
END PROCESS;


LED_1 <= SD_SLAVES(0) OR SD_SLAVES(0);


SYNTHESIZED_WIRE_575 <= NOT(OUT_pDBIN);



PROCESS(SYNTHESIZED_WIRE_565,SYNTHESIZED_WIRE_724,SYNTHESIZED_WIRE_725)
BEGIN
IF (SYNTHESIZED_WIRE_724 = '0') THEN
	DFF_inst512 <= '0';
ELSIF (SYNTHESIZED_WIRE_725 = '0') THEN
	DFF_inst512 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_565)) THEN
	DFF_inst512 <= SYNTHESIZED_WIRE_725;
END IF;
END PROCESS;


ROM_ADDRESS(13) <= ROM_A13 OR ROM_A13;


PROCESS(SYNTHESIZED_WIRE_568,IN_BOARD_RESET-,SYNTHESIZED_WIRE_569)
BEGIN
IF (IN_BOARD_RESET- = '0') THEN
	ROM_A13 <= '0';
ELSIF (SYNTHESIZED_WIRE_569 = '0') THEN
	ROM_A13 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_568)) THEN
	ROM_A13 <= Z80_LOCAL_D0(2);
END IF;
END PROCESS;




PROCESS(LOCAL_SD_SPI_CLK,SYNTHESIZED_WIRE_724,SYNTHESIZED_WIRE_725)
BEGIN
IF (SYNTHESIZED_WIRE_724 = '0') THEN
	SD_READ <= '0';
ELSIF (SYNTHESIZED_WIRE_725 = '0') THEN
	SD_READ <= '1';
ELSIF (RISING_EDGE(LOCAL_SD_SPI_CLK)) THEN
	SD_READ <= DFF_inst512;
END IF;
END PROCESS;


SD_CARD_CLK_DIV <= NOT(SYNTHESIZED_WIRE_726);




USB_DATA_IN- <= NOT(USB_DATA_IN);



SD_CARD_ADDRESS <= NOT(SYNTHESIZED_WIRE_726);



SYNTHESIZED_WIRE_574 <= NOT(SD_CARD_BUSY);



SYNTHESIZED_WIRE_724 <= SYNTHESIZED_WIRE_574 AND IN_BOARD_RESET-;


SYNTHESIZED_WIRE_486 <= NOT(PORT_SELECT_6F- OR OUT_pWR-);


SYNTHESIZED_WIRE_565 <= NOT(PORT_SELECT_6F- OR SYNTHESIZED_WIRE_575);


SYNTHESIZED_WIRE_559 <= NOT(SD_CARD_BUSY);



SYNTHESIZED_WIRE_576 <= NOT(OUT_sOUT);



SYNTHESIZED_WIRE_90 <= SD_CARD_READ_DATA- AND USB_STATUS_IN- AND USB_DATA_IN-;


SYNTHESIZED_WIRE_568 <= NOT(SYNTHESIZED_WIRE_576 OR OUT_pWR- OR PORT_7-);


SYNTHESIZED_WIRE_677 <= ROM_A13 OR ROM_A12;


b2v_inst53 : 74157_37
PORT MAP(A1 => SYNTHESIZED_WIRE_577,
		 B1 => SYNTHESIZED_WIRE_727,
		 SEL => SYNTHESIZED_WIRE_640,
		 B2 => SYNTHESIZED_WIRE_727,
		 A3 => SYNTHESIZED_WIRE_581,
		 B3 => SYNTHESIZED_WIRE_727,
		 A2 => SYNTHESIZED_WIRE_583,
		 B4 => SYNTHESIZED_WIRE_727,
		 GN => SYNTHESIZED_WIRE_727,
		 A4 => SYNTHESIZED_WIRE_586,
		 Y2 => S100_A9,
		 Y1 => S100_A8,
		 Y4 => S100_A11,
		 Y3 => S100_A10);


SYNTHESIZED_WIRE_91 <= BAR_IN_ENABLE- AND SYNTHESIZED_WIRE_587 AND SYNTHESIZED_WIRE_588;


SYNTHESIZED_WIRE_587 <= NOT(PS2_STATUS_IN);



SYNTHESIZED_WIRE_588 <= NOT(PS2_DATA_IN);




IO_OUTPUT <= Z80_WR AND Z80_IORQ;


IO_INPUT <= Z80_IORQ AND Z80_RD;


MEM_READ <= Z80_RD AND Z80_MREQ;


SYNTHESIZED_WIRE_728 <= Z80_MREQ AND Z80_RFSH-;


b2v_inst59 : 74373_38
PORT MAP(D1 => SYNTHESIZED_WIRE_589,
		 D3 => IO_INPUT,
		 D6 => Z80_M1,
		 D7 => Z80_INTA,
		 D2 => IO_OUTPUT,
		 G => ADDRESS_LATCH,
		 D4 => MEM_READ,
		 D5 => SYNTHESIZED_WIRE_590,
		 OEN => SYNTHESIZED_WIRE_591,
		 Q3 => OUT_sINP,
		 Q6 => OUT_sM1,
		 Q7 => OUT_sINTA,
		 Q2 => OUT_sOUT,
		 Q4 => OUT_sMEMR,
		 Q5 => OUT_sWO-,
		 Q1 => OUT_sHLTA);


IOBYTE_OE- <= IOBYTE- OR SYNTHESIZED_WIRE_642;


SYNTHESIZED_WIRE_595 <= NOT(Z80_RD- AND SYNTHESIZED_WIRE_728);


SYNTHESIZED_WIRE_672 <= NOT(Z80_IORQ AND Z80_M1);


SYNTHESIZED_WIRE_667 <= NOT(OUT_pDBIN);



MEM_WRITE <= Z80_WR AND Z80_MREQ;



Z80_INTA <= NOT(SYNTHESIZED_WIRE_672);



OUT_CPU_CLK- <= NOT(OUT_CPU_CLK);




WRITE <= NOT(Z80_WR- AND SYNTHESIZED_WIRE_595);


SYNTHESIZED_WIRE_590 <= NOT(WRITE);



b2v_inst7 : vga80x40
PORT MAP(reset => IN_BOARD_RESET,
		 clk25MHz => 25Mhz,
		 FONT_D => FONT_D,
		 ocrx => ocrx,
		 ocry => ocry,
		 octl => CTL,
		 TEXT_D => RAM_TEXT_D,
		 R => VGA_R,
		 G => VGA_G,
		 B => VGA_B,
		 hsync => HSync,
		 vsync => VSync,
		 cursor_x => CURSOR_X(6 DOWNTO 0),
		 cursor_y => CURSOR_Y(5 DOWNTO 0),
		 FONT_A => FONT_A,
		 TEXT_A => TEXT_A);


START_SYNC <= NOT(Z80_INTA OR SYNTHESIZED_WIRE_728 OR DFF_inst92);


b2v_inst71 : 74244_39
PORT MAP(1A2 => pSYNC_RAW,
		 1A4 => SYNTHESIZED_WIRE_729,
		 1A1 => DFF_inst97,
		 1A3 => ADDRESS_LATCH,
		 1GN => SYNTHESIZED_WIRE_598,
		 2A3 => SYNTHESIZED_WIRE_599,
		 2GN => SYNTHESIZED_WIRE_600,
		 2A1 => OUT_CPU_CLK,
		 2A4 => FPGA_IN_INT-,
		 2A2 => 2mHz,
		 1Y2 => FPGA_OUT_pSYNC,
		 1Y4 => OUT_pWR-,
		 2Y1 => FPGA_OUT_PHI,
		 1Y1 => OUT_pDBIN,
		 2Y3 => OUT_MWRT,
		 2Y4 => S100_INT-,
		 1Y3 => FPGA_OUT_pSTVAL-,
		 2Y2 => FPGA_OUT_2mHz_CLOCK);


SYNTHESIZED_WIRE_613 <= NOT(START_SYNC);



JMP_ENABLE <= NOT(JMP_ENABLE-);



OUT_RAM_WRITE- <= NOT(MEM_WRITE AND SYNTHESIZED_WIRE_722);




SYNTHESIZED_WIRE_668 <= PORT_C0H- OR SYNTHESIZED_WIRE_667;


SYNTHESIZED_WIRE_32 <= NOT(SYNTHESIZED_WIRE_603);



PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(7) <= SYNTHESIZED_WIRE_604(7);
ELSE
	Z80_LOCAL_DI(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(6) <= SYNTHESIZED_WIRE_604(6);
ELSE
	Z80_LOCAL_DI(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(5) <= SYNTHESIZED_WIRE_604(5);
ELSE
	Z80_LOCAL_DI(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(4) <= SYNTHESIZED_WIRE_604(4);
ELSE
	Z80_LOCAL_DI(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(3) <= SYNTHESIZED_WIRE_604(3);
ELSE
	Z80_LOCAL_DI(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(2) <= SYNTHESIZED_WIRE_604(2);
ELSE
	Z80_LOCAL_DI(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(1) <= SYNTHESIZED_WIRE_604(1);
ELSE
	Z80_LOCAL_DI(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_604,ROM_OE)
BEGIN
if (ROM_OE = '1') THEN
	Z80_LOCAL_DI(0) <= SYNTHESIZED_WIRE_604(0);
ELSE
	Z80_LOCAL_DI(0) <= 'Z';
END IF;
END PROCESS;


b2v_inst8 : uart
GENERIC MAP(CLOCK_DIVIDE => 1303,
			FLAG_HIGH => 1,
			FLAG_LOW => 0,
			RX_CHECK_START => 1,
			RX_CHECK_STOP => 3,
			RX_DELAY_RESTART => 4,
			RX_ERROR => 5,
			RX_IDLE => 0,
			RX_READ_BITS => 2,
			RX_RECEIVED => 6,
			TX_DELAY_RESTART => 2,
			TX_IDLE => 0,
			TX_SENDING => 1
			)
PORT MAP(clk => 50mHz,
		 rst => SYNTHESIZED_WIRE_605,
		 rx => DATA_FROM_USB_PORT,
		 transmit => SYNTHESIZED_WIRE_606,
		 data_read => USB_DATA_IN,
		 tx_byte => USB_DATA_OUT_BUS,
		 tx => SERIAL_DATA_TO_USB_PORT,
		 received => UART_Byte_Recieved,
		 is_receiving => UART_Busy_Recieving,
		 is_transmitting => UART_Busy_Transmitting,
		 recv_error => UART_Error,
		 data_ready => UART_DATA_READY,
		 rx_byte => USB_DATA_IN_BUS);


END_SYNC <= NOT(DFF_inst95);



SYNTHESIZED_WIRE_729 <= NOT(Z80_WR AND END_SYNC);



SYNTHESIZED_WIRE_599 <= NOT(SYNTHESIZED_WIRE_729 OR IO_OUTPUT);


SYNTHESIZED_WIRE_600 <= NOT(SYNTHESIZED_WIRE_683);



SYNTHESIZED_WIRE_603 <= NOT(ADDRESS_LATCH);



SYNTHESIZED_WIRE_598 <= NOT(IN_CDSB-);



FPGA_OUT_CTL_OE- <= NOT(IN_CDSB-);



FPGA_OUT_STATUS_OE- <= NOT(IN_SDSB-);




FPGA_OUT_LOW_ROM_LED- <= SYNTHESIZED_WIRE_677 OR DISABLE_ALL_ROM;




PROCESS(OUT_CPU_CLK,Z80_IORQ,SYNTHESIZED_WIRE_609)
BEGIN
IF (Z80_IORQ = '0') THEN
	DFF_inst92 <= '0';
ELSIF (SYNTHESIZED_WIRE_609 = '0') THEN
	DFF_inst92 <= '1';
ELSIF (RISING_EDGE(OUT_CPU_CLK)) THEN
	DFF_inst92 <= Z80_IORQ;
END IF;
END PROCESS;


PROCESS(OUT_CPU_CLK,SYNTHESIZED_WIRE_730,IN_BOARD_RESET-)
BEGIN
IF (SYNTHESIZED_WIRE_730 = '0') THEN
	SYNTHESIZED_WIRE_683 <= '0';
ELSIF (IN_BOARD_RESET- = '0') THEN
	SYNTHESIZED_WIRE_683 <= '1';
ELSIF (RISING_EDGE(OUT_CPU_CLK)) THEN
	SYNTHESIZED_WIRE_683 <= SYNTHESIZED_WIRE_730;
END IF;
END PROCESS;



PROCESS(OUT_CPU_CLK,SYNTHESIZED_WIRE_612,SYNTHESIZED_WIRE_613)
BEGIN
IF (SYNTHESIZED_WIRE_612 = '0') THEN
	DFF_inst95 <= '0';
ELSIF (SYNTHESIZED_WIRE_613 = '0') THEN
	DFF_inst95 <= '1';
ELSIF (RISING_EDGE(OUT_CPU_CLK)) THEN
	DFF_inst95 <= START_SYNC;
END IF;
END PROCESS;



PROCESS(SYNTHESIZED_WIRE_615,SYNTHESIZED_WIRE_731,SYNTHESIZED_WIRE_617)
BEGIN
IF (SYNTHESIZED_WIRE_731 = '0') THEN
	DFF_inst97 <= '0';
ELSIF (SYNTHESIZED_WIRE_617 = '0') THEN
	DFF_inst97 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_615)) THEN
	DFF_inst97 <= SYNTHESIZED_WIRE_731;
END IF;
END PROCESS;



FPGA_OUT_RAM_OE- <= OUT_RAM_READ- AND OUT_RAM_WRITE-;

FPGA_OUT_A1 <= S100_A1;
IN_BOARD_RESET- <= FPGA_IN_BOARD_RESET-;
DIP_7 <= DIP0;
IN_SDSB- <= FPGA_IN_SDSB-;
IN_CDSB- <= FPGA_IN_CDSB-;
50mHz <= CLK_50;
DATA_FROM_USB_PORT <= USB_RX;
DIP_5 <= DIP2;
DIP_6 <= DIP1;
FPGA_OUT_A2 <= S100_A2;
FPGA_OUT_A3 <= S100_A3;
FPGA_OUT_A4 <= S100_A4;
FPGA_OUT_A5 <= S100_A5;
FPGA_OUT_A6 <= S100_A6;
FPGA_OUT_A7 <= S100_A7;
FPGA_OUT_A16 <= S100_A16;
FPGA_OUT_A17 <= S100_A17;
FPGA_OUT_A18 <= S100_A18;
FPGA_OUT_A19 <= S100_A19;
FPGA_OUT_CPU_CLK <= OUT_CPU_CLK-;
FPGA_OUT_sINTA <= OUT_sINTA;
FPGA_OUT_sM1 <= OUT_sM1;
FPGA_OUT_sWO- <= OUT_sWO-;
FPGA_OUT_sMEMR <= OUT_sMEMR;
FPGA_OUT_sINP <= OUT_sINP;
FPGA_OUT_sOUT <= OUT_sOUT;
FPGA_OUT_sHLTA <= OUT_sHLTA;
FPGA_OUT_pDBIN <= OUT_pDBIN;
FPGA_OUT_pWR- <= OUT_pWR-;
FPGA_OUT_MWRT <= OUT_MWRT;
FPGA_OUT_RAM_WR- <= OUT_RAM_WRITE-;
FPGA_OUT_DO0 <= DATA_OUT_D0;
FPGA_OUT_DO1 <= DATA_OUT_D1;
FPGA_OUT_DO2 <= DATA_OUT_D2;
FPGA_OUT_DO3 <= DATA_OUT_D3;
FPGA_OUT_DO4 <= DATA_OUT_D4;
FPGA_OUT_DO5 <= DATA_OUT_D5;
FPGA_OUT_DO6 <= DATA_OUT_D6;
FPGA_OUT_DO7 <= DATA_OUT_D7;
FPGA_OUT_A0 <= S100_A0;
FPGA_OUT_A8 <= S100_A8;
FPGA_OUT_A9 <= S100_A9;
FPGA_OUT_A11 <= S100_A11;
FPGA_OUT_A10 <= S100_A10;
FPGA_OUT_A12 <= S100_A12;
FPGA_OUT_A13 <= S100_A13;
FPGA_OUT_A14 <= S100_A14;
FPGA_OUT_A15 <= S100_A15;
USB_TX <= SERIAL_DATA_TO_USB_PORT;
RTC_SPI_CLK <= SPI_MASTER_CLK;
DIAG_LED <= SPI_SD_CLK_SPEED;
FPGA_OUT_SPARE1 <= LOCAL_SD_SPI_CLK;

END bdf_type;